`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KjBO0tzHYKmFz+A6rqum84g+M5WFU0kFm4+9K8LdlsLYzV0nngEL4jep524QSuXSoSvZyB9EUMwc
kTLH5ij1pw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
edJqp/g900AsxfZU2BonoTWahObkFSINUtQ27mA19DFwQgOzeKWKReLqpKmVUqGeZPvfHC9/kaKP
tKQcjwtRT8veKjMbit3dubyXZrylnJZlMF68gkZsNKIFGCsJmH5O//nXHmBxeIcX1VAKR8Kr9bzb
9kr0dXKII8B7kkypmzE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
prrmYtH0mJsOZvaKbY12+aE82amXdifq/PlZhaKoSzNg9RAatFfMv7wDlt/fpLNtv9Qey7tbMUl8
MkDCxdbH+Rwcuw9sPCvyLMoIiUOAIuIeJrdLqqd1RbvedqMyDzRwwAnGOASLWmnlguCWzS2Pnwvz
vGnbtuhDQTnW885p44jjGwH+MlD3UjnmN6CykUPvxFZ7FcszS4WDhWNmpeU9LlxdsauS1Vyo+gFw
dajhEELJZAapvwZezOLsB6feUnatwWO9pIMPcuNpptKclbsp0+TZ2ROuJSLXF43lqIbjOCraKj/8
mHdQf7oU45lg/R0U4r49d8BbgiC4QUMXbm+tiA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
34obdx+3WX6Rhrd9YL0JFfGkdbdojfRJDEPdW0F3Bzwx0aCtsjTdFFmk6CbLjcBqkXZ5kVy3bitG
rkvVRX1d+lPY/2+8PXXoT0o0YpuNnDJMqJt+Xf2iJXQCsFP9O72dJrOGd91dLvEPOV+THlGs70r1
CelnPAGIWlubtMMOZUo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oE480r4SQjTvFUus7cCDxBRnypFQ6MKCoEgb64GS7nGOqBgyV1LfA9vPQiVjLMOST35nGj0/ddYR
Ta4Z5X4pv+g7OyjJKH7xVhZVw+61bRvj7bDTydwIqgcbS79OoXN0TTdu80hawRESaD+O4cgSYjut
ALGVTde4Cp43wt2hLAT/bFPswr/eg0WAz/HjBD++Qmm4YsMHgONAfiju0DQlW7fpeymHCO1Ucb9l
eF7FW/G/eecgeJtWYVFj31mkp8SqVP3D9Ehn29JKNJiUCBNy1/QohdeydCjuKIKSiEyunFLfh/KE
M9k+4O21klg75W/snJBQbtyW/SAh07cdxEPcbA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GSEQ+2k94SIzE8jZjjqbUn6zyZIVVMMPEXurn3kNUQzj9WZDEimOrNj9B2Y6rDGB5BYSCwrhIRaN
TXlaMBSuD6q16zpjPsERo72vwghPswLGmq8Ffa0BgTi/w3fStsI0TGJGtmWG4CejBXcIA5dbVdPt
DwwS0V18GxyX5P+UHGftIj+lhSH99agN6FoYNq7SiFqqze6UZv4zRHmwGSduFeiz7q4qvSd/+1fk
nOYi+qUnIcESfQGzoqIycVnspHzkQK1D2JFDedglr2VHstfkd7CeLLyIAZH6oom1FXiubsrGX57h
lJeyCfY2lEYMfqt9MPl2wormDmNt42dS7z+pKA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18704)
`protect data_block
hQ3CT7HOkkrGdFbh0TSqSIOeIzQ/cJlSOY1X493Pc9zXawjFwigWvC1Q7S5esKr1zAGkfEuKCKkg
ZAWjFI+twdvhxMB1ilTSn5P07vAOsLQqrhL5Mzd//qspzYfac5Ys14iIKuNhIFKmBJ4qyUXL65ct
KyXGXjO+thtKBnReZcys6/7dZ6vsS7ZXUicU9Ppg+MHwGHcScj6Hfyko5JisbxNB+6sKye98VxAB
4T0y7wGWl8W2A+tdJBe3ddTO9x5V/YTchkjwwuiFQRJqeYB8CgtkTcVHcF6rxJd7epTgVKuW19LE
paeWG7Q/OG+8O9jQgEPqxD5wzTD/RB0tGzribx98ZjCrUNUvg0IibWN1i1S72SlFKXdb8qsfr2vz
nBqwChHyjU7tth+rB/Jow1QCdj9R5LQaHBnMiWXJGs7nSUMEx2EdsvL/Xl0j2VC2e0AmUpwgQ/YM
VMA18slyVR+7JL1s9AtsHxNHCXuhBO9w/AK7Vl9i4Ywj2vUamPNwk00DDwyQYYRHLzkv+D3vX9fF
oF0pqDWEO6Gpj/aCkwaGO0ISZcBxRGruUVMreCcPMssp/VkxhCGFf1yxiZHS8b9ZyK3F3gvJYLwJ
db6VqWrBP+ORK+bBKCs1yPnVWYs5t7grbHdLu+fBsFyyPL+IiOjzUqKz1tdqsQ1RSnyIQu5ZsU17
Q5mTgcE9GHikzQ8xCi+Mxv1p2Wi6Qau9TzyLfVbr41CSgd0VtRkRT42jURNNs/2qrYEOefDplnn2
ZOyeYRlZBpD5v4YdAVqWg2Wo4n9t2kfLhycJDSeRy+DOQCFdb+WAmzyWtI4AIbwqwYE0NApVaKfd
vd4Omnk31JvoGxzll3tptT2pcDbO2dWZkx0oOkRWIp5mo5NJA0LOCOj2zih4DBe8ciK0zRq7EoYA
hls0ZSE3b1Cn6Dg62g6Xz2t4q9ybdZue/LNejFxxu7cNZ56bc5Lx1FtXx53o/DbB297luQBWCHwU
KaWaAIok5GRH/l+xQ+WsITJvPxvyFqs/+VjNUWYQty06+wU7vs+dTsB7ocWWHVz2/XQSXd+t9Hsr
6NVJlNfS608KQj3/hRPzf/i10bu0nYzyUrdPkM/yAOOwy3w8y5qtk2v2nkE7RR5R88FROblmmFk+
negrLTeHSU12YL4eXxzmjWTHgsMk8NOAQbspVbQ7yQDq9V4VCDUQQeUt28IUk5hge8pqNLwTZVg5
HgIXQAJ7hV3C/YdIHGjl8W0wwEIH9qBvJ6b6DtKt7lDf9KRYyXhVStwzoZarwSzba5mYO4H0IJ15
g9QEcef9RAyLLdvJfQ+gxyfxJwJln2t8RsW1Dsoe0QTvKCua4HsyBVmNzPppL+pyms9lDqa2HFCg
8r/jnMc7QXMbi25pJWrx8S1JjZVHYef1fJVKHEmKX/Rmn7+xP+nwDicBsmMmXNaPvIzp7Aqrm5ck
Ju42BqmssNUHluC3X1IMElql2MiPOfT0GOMBYIw2X4uo+gAoASrEBDGKQEQoK+meqeIuQIOGVLLo
QjEFns/Apk9Jy+I683mqpg/ghLKAPe7i2WQEMs0/3y6LgFuBMGmSP828ZbfMVVPkceF1aHLO8FEs
Hxx77Rr2aL8BRdg9oCDMFnUF5g3KQh2exZgops24DWjhO/JCFTuqspIQhUn9jvjUbliwtVeIha7a
9adeavFjXw7slNyBDaYMSIHoXidyuXuRqY3KbBKzDjTBWMe6IDFg6f6Ixv/8m5YpNsac7tteFwNE
jtvn1LKg9vjkoUh9XFb7j+C+WccksJ9hF6icKZf2HfkJqAyIx4PHIpWjHAqfZxe5NZ14sL4/dl63
viPP+zgw9PTEwTPj7BFyHtTv/YvjSwtH0cYZtXfr0YXSKJeAzOggNDo5iY/T53MjK0djMY8l8mOu
JW0M1HuyhNTxwYxness4AEoifyuXAZdQXr/3qKdq1CUhqtUDtMaF3NWBlWqo41I1LFtgmmBlHuLb
c+K1FLCKqZGxKPRwyxGv4AL74he82ESXrsi7BjA8HlyAlncB0Te0wcYO87ZElDuj6dNPGom3gi16
7x0Xtk4vhmBAemwxZ7AocOrtgA91VJDknAKcY07HQy4QPSs3WOa2WbCc8ppniHcDbtbkXTncbtGL
pWe6dAvMcIsYwjFx72GAImHZ1jIrYmzVq4UWGGMgJm1bPRV5PhNnpZjhd1BWlOkM4Pm3kXs2QBJ/
jqO9n8qUT40F2z4MnC7/qG1GcH4jFrIV8ypWMZqOx8kxG8ZWTrFAOXg8yO5psPvFz1Sf1tzTUquP
aVey5flIiy/4npq3G9RFiIIwI8RQiFvlQ7ClCiDNfcg0jMPYNWKE8svuU8JNF/dczGpbwn4zu4bO
O4+6wOimwYD8oz7CC118VWgu+oET+Dn5YtZmbAP1UhWVMQQ0HpxDwsJokjNldhLNq82oYsNgQd+q
V88YayfiY6888aqr7r7zOW+pDaWGA0A1ciUSCe9dSdF+SSy56yImln+SjkP/Rrrur6FoDGx69ESM
0aUNFx44nfwUXuy/84dAazMrLNCJlXK0EgwR90qvBLEM+VjY0PeJ3aph8ekO7HGo/rhZAqEeZbr7
axg7OZdIABm+PQYEjbnM6qvWxpTAWPe6ubYOWxXJ3FS2vw/tzN4VqhGCRVfdGtvDyLtQSU2NPAQJ
sZOOa5R+JRUPEXq+l/yxbRJSPgojwEmaEORxksa5cekJ0uGph1u98rzDiN1fdC92nvtN+0aqowGq
AIn+6TrlgdGbdt0nHEOIB5NzNu7qG79ZCnCkc2QqDMB29kGKf8y5Pl6xLxcib45Qio2Jc5vM0FcS
xCAbUFVy3wipN8CZnA88Lcx/Kzt8FvbkKS0TsaElyfkDZxDVHVYoFGwl7VpmLq7ZXPTzgSX1UUKP
UQiuQpiMUJvexLVz9Jp3/tDbeCjsDwGR2LP5yzIMV9oqz1DIg/PuX6CMsVgJUkJipdh4hZ5HEuvs
5LbTr9PZDT5Fu/1VYqE9l32GEJfrYdeNkc0O+4kt0u8upAkPmgRwPcZqhhTNPWAgrj2T0+eiAOTy
ZVJCnjxlCnLsoqt46fLx1B8XU9JD2ld5CZeUvcd2AfXjkK2wFNxWIeJTbXKVZVYrz1GwaocVrhvB
sv2MZFrqStEAAukMLsjMlfY3HKtsgXjuMgktup73Q+uJXgUeLFGo+3Xm/nnhA+D4Xn8W99zzwPS1
D1Nl23lXLxM5CXNIyZZKT+CJUoT0Pde5RQ/mGXegrMltGXRAHChnWzONOZrTk/5F5IWVVCmg1eq4
eSbjU6O7KrDZAtWhWmwkW4fwYHrc2dojAIqXK66f0eBSBisNp3G+xHYvj82B/DHUyZ4Nl6SQ5Vg9
woa2YjgyPMXLfC5oDVe9wMsnAFSlLo5XMcQX6twgvq07mj94RVPbX9Pk2mgyjZZiFApsZUgnVHh8
5Hw/15rzuzqYEri7XWSM01kMWzZrKXLyqx1sR5FTVpzxrTNpDE94k6D+3sePmz9EcQIenGGM2mLy
//LNoocMmpOBzm+ovyYnDxNNCnwLmhEX1v65M05YP4YrxhCJwr9aTa/hJ/KPc2MmV/hHu/0fNb6f
xAP1D8WpGHY5Wi7o4l1c0ug1i1RYSNYDdzDqYkDjiULEy5fUOs2aEM+6xy0/0m+bXMoH++A6v5a7
veErnbULtoFz1RTQcUIKb1AKRsa+o2n5KBbY+H0yMzz9zNJovlj7zNBnTgt3DNsgSclhWWVWYpjL
Jy/Xh7vRTSLEmL0I/FQCkZ7hFLEy1ixVSB2ySQfOg1stuxjojDiaUDdHNeNW9Nv4lbJyqKaDqWYg
4XEcEElHFyLBnn+W9ax/zR4pM+XWbHG7l04RimR1a8xw50CbpSIWu2LbqBuCLIwoaYC3lJz30s/B
vHjbfk/TMdeahK8uBmrVoaqfauVgQjTxeDO1M2fYk0PY5ZL0p/9aGCKQ8n/rowFLjGG6fyzGSpbc
NDlTMt3NVY8VvnDNdShOsCF8MXoL8q9stfz1yuv62zL8ccMzJwk0sxO7JrS34e65C0n04KSxCjfs
k0kKAicjRrgEaE9UUIq5vOC7Xfkl0jmOaKZk0Dq3kE8ZHMzr787z0xrQzdhT55KP0VO6mG3yEHjl
GNhLx97pAE3zXzHGYYFS4eDCJ+pZ23J+Gxu7DufD6bKuNw0v4w7Nfutd0Hnu5DG70U4tsCOuIeQa
Sy0dWsswxM1oRdmqPx6tjmOpuCeD/eK6PEcCux+1z8jzw8rf1DP6OXpxiAwUS0gieyesaOnnVFFa
FNO8I2LlL3O9rC6E9Be6NwwML/zOocpmsV7X52mqVZV7l3J5wCAshOJbAYK8pAFFdvdG496t5bey
h+mnw8o4IprexAuzmoU1LrR8QAgyPBZ/+HGsMHbBe1gqnrbGu5lPoAcBiWAv80nQ3gk+bw8eEaRR
RzSylH4etS49Pwu6ey2/WYN+k1o2YJmx2cJCOlgT0IXxI9eAxbG6cBBKnSMkVDPWRjalm4IYxVfm
dJbFvqYn1BYaupVFVmbFegRBQtG+Cm3kdOacj4oIlky6stB7+QYYSOZlHcHztSX6d4Hemu6Lo+LV
kvNgoD0VHXerZ7M1NLfwniOWHT6Oy3NK+i1eeFBEZH/ZgVDd8lnHUd2Mtxnk00wz50RyRmncmTbL
p0UkTc6Q+RmmXj1nW3UBFRS6uDFCI628QDQI3y0VfkZwzcb9MOKEjx3LnXh1lg0LYd/mAdbbbnBS
jwL06aS0VoAXuDfq/CF2hp46wfC1dF96OAdVIGvz1dhPpJkdVxlGl+6DzW6J487qwdfhqM0vWSe8
QujgfA+ICkSWbBuiNW0xBrFQA4erH3dyhyhP3EEPntHHzEJANJ10lw1XfWhj/QYLX+GqAUkNZxVp
iPNkPSUMc76PVIv/+4Ig9lOso/spmC8PgGfLM3fPDVXA2DVXe3Va49dbbkpU/Idp5C0SDKleOElW
FTMbdvVhYMpspsyI6rPv/w7EqD5f/J89au3soEuCeHsH0nBqaRC8wC7RH7+DmTejIGa+/NY6g+ZY
EvsNROqwJh0bnLslflmBV8l5kt3m4XTsy13wXVxGmGUs5EBQtRuGRl9gRi4/ZazT9Uesen3qPqdj
fDQrKzUdiV2GCEn/R84Cn19JM4P4V+k/9zhakzm6QsMaGKJ9hdGx5eJ6mKUw5TktN46sy6doVk5A
6pwufKgaSNvWvygr7rnpNphlSTGdU/EAAw01VyxoPWtp7DzfNO+mn/ylDUol1jUl9RXItGSSnJDt
cnj1jhnd2nOWedUfKMMHyTideGb+l/iN6DQS/hGoFk7RwlRsS66Z08fLuXGddbDya/SW+sudGo/+
PGaUBamoPpVcWyaDWzLyTI1CUkMbiRoNiIWQb7h8Lih+OQqcZSIHS521VGNFaunsr2ul9c+aUbkK
mCvEFKdyeFO9C4gYiRSJJmHowCEaJnOPtLrSto0QMvWagSH5J36x/bUBpfXnhU0NDZgXxmGK0DN3
O2zLTzngAtqxEa5XtlU3DkI6MdsOQOl25yLNo5s/Suc4yRS7q2HUDH76oqAyRTJw4JRsOlOkjI09
MReCyuCDneGkGOajzpoaYkIu2ai2UuiOIpHr/YaOXZ4CHd7/TT7c0/aqZLvfLsAfzV//PCFYvXRX
kHaaEUIhoakArtxckfrxTjt8mVE18nwf91n0lI6JagE/H3F6xjzor4WmGgzByVfYI+B6415TajQ7
vGft4IU4P0og2d30N0wtBam+6s9nmt6Xt3tGSbPKqmTc9qVnTwddC58kjBo5SqlsMuSdeUa+3sv2
YsBZVAPRcocamKs8/ruT1qyys7BXUk6RoOjWdWxMp0dT9jhyYQ0gFQ2sIth18MirtQBCzg5EzzPJ
uCo+fK2JWUBfrvcV2rcJNpIsPqSVG1rkjA4P0HrMvC5gbojNyDH9zQ8J6Cjf1epkN/74ZyUhSgsk
LaZE6Q6eXuFRYyHivXr+NFl/mezT9CkvRtysH6jjwNMqzsaoxh8WJ82zZ3Z83Iscdq3fDdeJflng
yoH8hXreupV08QMrMrjh7ZwwJHtBGAy8ep8ufbH/q532rfjg2/FjSwaQjdwQbdodKmmluc+lLPeR
w3NVzBxJR0JerP2ixKWaUOnHBpUH3whVw6OBKlXyNk+7Wy1tul1ZX0fblYqImF6TAi6LEl/HCABW
PRpJdTuv9rjxbLkQdA9bR/nEL8jQfi3GNxQzPnMLnGvETiCEg0FPXm9k0u7vdLIvF6DRbt6bwLVz
AYhBXYsjEk83kmw/jxPodsZRePjgCryQjx5pa6+OqQWvg5Vk03PqtMiJD4Lt2tgrt/Rav/jBefOp
HZafs+n0+KOqYRckWUuvkcIzlkpDTPiDOEZ0CpVwgAB8/dNjkpkcaS/nHRu9F9VhwtNJZV78w+yI
deD1XvHu3s1rK8vCv3JwqQSYZ0dNanzUQJTFJ/1YWOVpuZh6FeJytDSCWDaSeVjCapTgaCys4csf
5EJfTWj0QZA+ms1DFKUbiQJr8C2UC+IG9mPRQpOVM9ktBYiNBhm2Bkx5f/1aMW16l8r7MVzac+t1
0yZhPjjmCoYhOni8eymWNUKmVHqjn+THXdyhb2LkSB0WozhjZuor2XLJSUManq/RXhm87YzIW2/B
8KNE1sVXmR5WPJO5h4L5eCyc9fuShPoZg5P0Me5a5tnM8im2udnrgOOMqH3V13l1zYSel0WmvQ9p
lJ/TUqh2CE6afvF8tQQqQItQEwAq+f5GCmSghdpJhq84aam2/sZ2w66JSkJHXWubRFNiF0jkSGkg
2/7Tygs4EgVSqxpIB1nbjr0GRY8y/ohzkNKGZTB+WVHHfPLw12juZE/P2fwTHr5nONt0aqFp0K3Z
+RX+XW57wnlTSZYtvuT7oHihv9gb2HmmL6yttdvMhJ07ThF+dgUcPFKG1nZukerh4QTqbtdNhO/a
0uhK05UXazZN7tVlPpBdR/a8dcevCqXn0JyU2F5OjPDayYOeKUXn50g9EszrSdX0NqfCzOKy+RF7
a3rvFc/onHB+bta1We6RAbtQALaZWCN+qp8sa43IEwnyJTUMFBqXNENEB5ElJUTnwg6tPLDWvPnl
1kq7Ocp0FSHVEh2G0XIai2TWC7M8aguoqaMqWOQ1K7iXCQX6e3P/UPWdiAnxCAGSZwEeucjB2qVV
KCFVev1qXFnB1drC0XNKX3GEvwjlD2JeXIGvM5kPP8oFgsJv+RY+BD0Y7t2sdp+7etxJdg08w1fR
vCJt0MLgdFU/qtC07Ug/VmKTmWr1URcGnbW0NyYOLHBi0pT3IeS1D2LuwkqMpTAtNvanRI2iXZmF
DTsFipj//NqdfW/iQsMJnREwwYh0o7cznEIbvPHI/GEJ7zip+6s4PAoCV32cLSJqbIec3fxFqejS
1GDgyI3a85KgNRCFvoxPKU8q0o8+yT9zzlahWIM6aM3G5vMmAzTBTzSEFNGg53aqzKqj3uewkr3I
tgoCjjj8cspkqUT1JxqjQRoFOGbJovfDkWdFtXMY7aZSBs309UdUR2cBqNYf36zmzk88kOYmbXCy
IIdIYbm/h+wNxjoivxePuoK8U5wFMjkRmD463BL71V0L/u8DPX4apKzmfcZOZuUkZF1KSubsmQvd
r9sc+jgvOU96pCJIuYK5scrnlgPl/nzhHPCtURoAD7pRMRZ9NnsXvrO3l0XEraZxbKUsP03gEf37
X1lsiNJ4xxgLP0trN//p4cQPlIkFifeSdcWqt5TYrR7/C7/39swqjVfS4whN/5TbpSnq3OcZn626
WifCjReObkhQw6nk8/M2fQjb/5/92eqDogmWaI/aLboVe9QGtTnZC+nE3d7KIJhwjP1kzY8eH3qh
t/99e94xoTbITW95uvrca98+wotMx+5ahXqm+MmL+Lf1Pj9dDES787ZSLyPvoR/OrJX0vJUt6wT4
dcmZsWSC834GyuDnXPYWf6z8OWCMiAfjwC8dr0+AwU+9ZKLc3uXXGd7RzXsbkZk2LvUHHUqx8ub7
3Sd1VfPJtbXbZ0QmAuoEkYkXNfu6ct0lr4PJyhcmx/wFKgUbUJ09x0boaAyI3kB5+fJGdYo1KjDp
5AGLFEV+OqPCbqrZ/kn46EAOAZ6RVXjqqS1gwCw9vtG+qcPGbvl3fLozIxUXgkfUy+irnd+KeeN3
IW6qhrYJJmIAqYhjRPxwPBxj82kC8dfJV+hsM8ACosse/JvM9jrMbgsMrFOlwQ+yhkF3cmD8H0XC
YaEp4IoL59P6pVhbvInbQHX7yPHYdhsW8v9glMUEo1bOZmif4C1BmitqAqSPJybCFOJ2UkvyTFQb
mhc4Gg2VQ4hmzUPNT+1GrQEeWzQyDt9Q0dlwPZYIXoeB27f3Y1ZMlOrfpTxnWbCRAu1GVKVNIdm9
dnVJJkoWfOvpOn7FNJLY1uWsUtEfy7O+pVtlvBHcZPm4i5d3rZmjWWE3swNc1lepKnb0lX2QHyQK
C3p93vkPV5bn54KGMiuqxpvd2ptq6j2AXqWdLpZNnHzx6UH0V9NB1wGvyRKILiCq2COLGOli+dnc
Yn3PPiD4cUTOMWeHmsuvkOAFSuPRa7+HxRtgM2JSBtOyM3m9rh/qK09mBtg4b091/5MJlt93Cpf2
jYrg0B7rqFu/JKWQ35G/A1rp3nH46KI0pCYyj7q8u962i2iDKJ8RTK3L1i0gs5A/kBky15PCjoxq
qSl/ZlsHviCyjxrHEmLQYsuh+v0xE1QWIDn7HerayYy8jQvfy33Mj8dqW3AKCjDsSk2Q0PSVy93H
8pE+qhnCd5Y8+1X8814YptZQ3Ds1cIO8F9F6CPzPa7IY4gC4UluZrh70BPYMdyssxzNDDk2bpCX1
iH5bELGYax8SuRAn13KAMjZ7YYuJ0ZoC7UBrr3lMfSA4fZ6oNf3RxOkKV6uG0nVkycOy1HB2qg/i
2dRzmszc44Sg2YTumB0oq4BbmeaSZnR3ThYi4qq/8mCOwgZbVei1549oi6PVsvq920alAtG46Bwj
Ed88nhi35e0FkfIWs+TQnPUj+2myl+2TFnPygvCrQ7wRJ144JBh8Ok2xomSOAEXhG9YvR3uJ29Py
ea3mwtw9W6DNCdw8DFj8Kni/3IM3CtddCOIoGqrxJ5ZA2nIdOvzT8n+fEn7BleJtLSAZPLbTpy7q
eUbp4YvjR1Ld8PREbvPinCuRzTAajqverjVRdXNJ8vemx0ohfKS4M+JyqnRibk7aZ56k65DIRpZY
ShirJjUImhzWReP2D/7xw5MWEKqCEq3jg1pGKhtWg3KXrxv6B6Ngga9cuJidn+mWgHSyHy+UK4kk
akxa75w2KxKRbWVBerMwDwVtJhjrCyoByYY6LlyRNxQ+PQLY8qIdAu5uGS6O2W8SChF5IUjXPJHe
U1IE7VZ27qtslZuUoYM2C7nAGGsiO1YbbjG6XZv6+mdP38mFhwle9AAl1aHQAST5ecFpO6Lo1X8O
HAiiw0LR+cBxd6fcOxDUjB78DKZYtFv8IXeZWK38Q+jkDslNf8xZbO2qhD2uD2kwq43tBZVvs9J6
/JnzsG6IyZaOqCAEhvEd5EmpO7Fz4TGV/Wtm2EObtXZv9fGHCi6rj0NVoKYciTGdLbsSqwaeCqhL
9C8ySz2pmRdh4gP2AfeBdhZawlEcUr/5O+n0e+j8d1b3x5dctJi5oXJCIEhhYOxlrksssFouw8U6
DZIyFLeZT8fiEoZctkFlR6Op6BKWppQ4iWvo1zIbyVozG7+zH0RLFnWgufK9qYYvVU1LlHgUad0J
7AtL3hC7fD0Nohvd/b8NHzYjRl1SV5EOB3gulP9+LwaWzoLU/bqobqiHTle1trVba5jXfYcKG4JL
8Y8CImFD82x5NCro81Knh1MZDDdpLYq1rVZ7lbQjDj6EdpRY8SWwcMwJGZUxqRRLjvndAO42X7on
wcoNqsI5UoQcOjnjhSvqIpPR29yxlG2rmuHac3HlqI2c/ZYibOsHpIZxIWowRAyOmyxrIxkZas7R
SptDTP/SyMvULOvbfSAM4EV7wAYtJgRu5TFIs0puZchXo5zP1oW8mcMJTEvqhLmubSQ57uvnplvF
Ty+sh6MfDKEdQKcULYxgJuRZJrhYH86pkC9IBI3bb7cTZh32bjiwe8H981NR9VNL+bNN4xSiqKgU
At2t3BxyMTe4tCoz3MLsMIcMpvzGtW+nbuBnO4E0Mc3m5KrNzeE1njjGaCquyqIayxKINNmOpQtu
jrtDkFP0vNepBO16JHE5plQr4Jre4rautM2EfO+zmnXUQSCwPQHt8qguLWfNn71AINsDKxu2j7Sf
1ndqTnPS7X2DzYXRKpZ25of6FP8Ay7Li/zn88fDPh7BakU34FP2hSS6Z6vabIAk5LEo1JUoPtR9F
I7D9OXrxNM4nG9E0uOdF/AlcK+OkHxl5bP6BTCz9BfVwgSG2yhX2kKikGe+OYoC/nvKrAqFIQzJ8
OLW/IxqJC6c2YhVs+9qCLJ5YFvvKnS2QAmG+DR495bP0Pna6AWMuh/uvvDeRjSoj025ogywZRwhq
5tYCwaTTAiFjTZqlNRDLgXEO2J7RP9eNqRkWykXbe8OBd+10qDq+aQU/A0cQnVu318ECsLB2J2/8
sS8GmyJr0EVbMnjRfJkTKMHPLsux4kb/PbL83UQiye4xARV9+pbi/bX/RDTnunCmMosytkRD1wqL
wT4AoAoYM2iT1r0fK1gPAjM0MjdxMjzGcg6flE8Inwqh9xyucQXCpd2kOAJDq4x3hQBlt2bcSl6d
64Gz53wdZxJ4vhIcr5nNtJfYG8abOQNkC5YXuFlx1jtjlyXFIltqX+gw2L09ES7DaG+C00JNWDvb
SbYtDWBXFn1iQQsriSgih4Qn8Igm7k1ILq7zjHmIUL1mT8tXYAjNUfHd3ss/HJxPuhVv92OYzw03
pZeMQ07fzS+OtxH0OEbLutn4OT0ED1GyIQ+TBOhQGdJSeDWmJwR5/xfGwEjahAkQ/qGpQxX0m/fB
lgEF/nZ7JvVkXd5REZ88QyAvZERyY3FKLoDex+4kE7PW4shTcpfmVfYr9QkZLW2CFYKYyqeHrZ+C
cyTay4fTLUxdL5wc+xs2unz+tpksLEsfB0liN19B9QtdRlF0vkM7WeCdPyJtsTaL50+M7iyyB2DJ
xUSRznz+Hs8xBQm9nafiAnViKDQ047UWS93Sg2oUGlP+a3wb5arcIHns47DFlMQt4CVIp6yqDLdJ
CanWSUaolRcN0MEpa9pT2d+pD+D7JruuIBf5vaOTEwpnJAyq2HAFFyKHgHAdgjeKlz3Ey0hG/ac3
NhgHqQiVg1Fj+7fVks9fRZXVajkDeQM/ko2NTPV3MjV38wIDPu9tNgd4RnHwnkyzj8mxLH6I4bOf
39DiLRTs6YU/o+ZXgcAgmn4Q6uLw5+DoO/KZCEYQU2DYOOIvnNJJuEgIPLk1vJaLY+uKyOUkt1vH
7UvgblrqFnVp4f+PnuaeyYWmHPRGDWLzimm8TocmUpsLe9LXfo1PGUO3q6WhjqFUe7WyH2Mc3keL
4P+GjiBCyx9vZXRDkimRFjsuUD/0ur48pouVzlW9VMXoKqjfH5ynTOYluFB5Dq4ezpMinZsAY4n3
NmeoPkhofpdUSHCCuU2tHM9q5Rg5zVY84Ihe/bfit2RHNVQ6Rrk4NWXBlZh5cUCe19KHZTurM/e2
vZ6UABDI+PESL9Z5WiSaTWhy7m0N/dh+aDGYwqdQk2h1DJevPWyYly46BtSUh4qv1DFXn1zB5/hi
6akExLaI5gXmkpdMpXtUoEGj3nEwn9/YqCdEYeJRcbq9Inm+uIifgXbPJkzYObZtRsPXWuzpGkXa
9gBOmb39BOANM4lL7T9DwPYM/iWHlJbjDgEwbiueQjsUCcrWuTLUi/+eaHOnzAI0eGX9kxF51whN
gge7SF/dPyC4j34zAx93tNwH1y6QKTdz/nnGlFzBYulyknGnu4ExulnrXIVdNb3UbrEms3Czq7MF
n93d8/q6KXZR29GkJQCXx5oAeYxoDqdjC78vzifMh//AnYxpMurIY/AEYLrHdkBIWBymoqIddGTE
AeMaidZEoP4O9HX1N2EXnIac9uRc3LafVEW5jVaxCzoRg3TE+uoTRtejpnNs4MRgJo4xzqQlJpe/
Y09SQSUF5WD6KbQl9aH3p0s2lrrJWEH194SRrXLE6Mj8mtc4KGbYipJzKnD/K+DVqwTozH5AtYc0
j7ghaSYxkIgshKhgarI9exfEvA0x9YHhKF1FrzMSqcz06m1ZSszhgjLnK4uALW+hQfreqHZ3MTRT
ojdU8EfBMxyi5AkSDgxP5IO5HHJGw0J2wDAZ79QBGfav1K0ie0nChBNRkWqsMpexN+fyLEtnGJ9B
O7KW05ZFEavbBqWjLDAakB2gKQXFoquvgLA3N8MPHLuP7fDS7ZUJ8sDGza3guiO4IDPgCmUxmVDx
i7pssCnk7EWYYzklzMg+yFM5SJihiubcOXYndhG9fUNkSVwirpJH+OAppd/e16n4VabUXyfulExT
jeHjDzFHH382pRRvVwZI9EOUATWdrV1mlYh0GA2P0W4mAYkwk82J2rGMJlnWO1KNEiYeLQuAt9VR
4m8yqpNDJtoIkv6auBrIrG/1GAHM4MyjdbyPACQdIyNvpo9kBExQU+lTeClhTjhyY2U6T9qMAwmH
+NP90z7F1/3ciZR3P6F5yFZgFgQLtVZ3+nvtH6yri6rcoeuMPJFM9SzH3yuN7KrWHXImWGmBhzju
Bat0MsbuajN/Fjo9Gnu2NEOJraTRlzdlloLixwN5nKIbjGJFTI3lszUvgspxUBS//QUfqtLRPzrf
//5DrFUN9HmFC2YUHott2cSHKGfcFBYKrQ/NnoBAeV48+C/Ax+i0P/y+PG2HNu68sH0gmWCTHH3W
vBsLozhU4mzByqKSsWhwdfPNNIYT0TllX+fwL6Q9XCfCoMTqY/PM5FMqpjpL3h0aN5/r1QfZWtri
5SRoq0YoWcCLKq9an0aqBW1kCcqZ1MSPw6zl+Nxq5g75iPMKxgk5A1A3Y6YYTM9a2jfj90GNzJ+F
jiZxZUt7WKrPujyxf8LHnwpdq+2HtntxTlU9CB43fK8S/t42mDNFr704lk+iqVzwRKH7ICVxEd7t
XK/TpsVlCepZ4y6UfTgKc+M5H5Pl2XnZY0YNIdcNuI1f4bAGf37kHcbf325nolcsOu/KsZm7RCgs
vWIGQrXFM7ZnJrGVWzmKBDHVQ6rBaIHTejjJN4dYjj9PX0mlDDh3x3LzyPQDflgttygDvnGSRkO3
HZkqOc0sbNDDsYUK5bStI2QOgpBWyNzrur3qppOuYzwJ5opq9NAORbLL+bLnpy7BmYNUNJe01isS
PhzNwvCY95DBhf+0fuNzEOoypN8/QMOAc9B/UrtcDEQBjS8d3QymRInw8oWHcF3t7AEXAHsf6yKJ
HoR1j6o5PQO8jr9ws07QZSFASuhe/VudhHM8oqdJqpi73AXL2/6GyociuuoGrP8WiWusEwwzN8nb
o+s+bSasAOV3BUBeg+C2GKIliJJeQkEU07cicWNpvdH9JJWpwjdwSZWTsDAW4n9JPqusLkARCZu1
4q9peea7d6A++ghFqlibSNuwfuKXRarJimEc/cf1EJWp2OjjY0V6FQj9HrJQ3q8P6E4FiUKtpw7L
Xb+jd0PpOYA0CVZI4Kx96McX6vuNUadVPSxl65XMeHk3yCBx/zd2cbTWFR6OwsVrhYO3enDGNWPn
5IrSt69ahU0dOMj9G4CkwuGnFMvRgQMhSaAxNKl9YyChANGJl6rxm5fdYOcubFwWK127tI5fE4ax
gu7JZs7qy3IO0//HSAQk1eJhPpnPqrpg+Wc6U0bFBSCUnQiW1anpqtFB4daJYUkJW8KuoqvvDQC4
csGfdC+wdAeE8UGjrvVbp/RLRQAaY6kiInFAJ3xf5FkK6fugBZrGHkEcLNZlNXzWoQyA1EKaXfdz
ed6/7pVCpDsxo6CMh/HLxXX7RXvhCSiyc3OcJEbpSjuuO1xsjEAzDFQ37Kl4MB7pvTm4xVVbYaeu
3wsFOy5u3OLWGThCfcUAQsSDhXa7fPiz1WSfR3m91BW9Ao+xavP7mv5CJhlYVtGfvoYe84Bb3/Oi
x2ykoG8hs3ssMQT4C/wh9jy+ijaYbbWf+3794G6fyVsSIBAL+CTdrlcOuZj4NzJNOsY+Rh9j9b/D
Woodm8Yz4NJ8hbfh6m6WWxI/OudaktnxwHWNtjMx9AGZF9gdaOEVluEt7eim3Z4dEGW1+CueKG+P
C41fdDYfoJqDK5mKoJIvqN4m3iEtRv4rhY8Zz8Y9rlbte5bU4+pwS56QbxatlVjQdgglfs0FRUqJ
cLVzcrJ8hutYvRFKbUyzd0NzQs6AA//TesxePCPr45muA5HcFAm4MtfalMfOd2wI23mDJKZDrTsp
9scQczdEBh3pmzmeK1WiJRZ7n/33tR+kA8fAPXwcZ1RuAbYEK5qysc+GNcZdW/pnH/nt8kIsuIZ+
0eiw22M7ToWUrHRajwVjv81BHdHeSTOFrPynoWA8MSzmYosNLyFgYm7YM6HNk9l8UlZkTnc6KbP4
YmMaaTzKVM7p0bDK9qgyBco7ffZuAfYSyvkmYik+wzMz40CoKt0YD2T/9vNyGi351INifEZng+tO
IJ73pl/4aUVnAj3bvmzrqYj/hpBhK1c7Uh4nuYV2SAjv7OziIIFWsbSCo7EVgMKOpkV9ueBlTkZf
/5cdprgzv2Ww9Q06XdD1cgHIei84RUALqg1M9RQFyYdTA2rxj3EfglbcSjeaCakZcHndjDKpFwZt
9WBnsw/dz6pqfEtz0ANGSSWky3GV5yWhIsP8SgtJW54oFp5+/UsY45HynT17JdGkaZ4O8JD0rY9K
AvdlZIom15Qx/mo+nilLDlzzi8XHyu8oFRKFMFGudgv9tUMHSKbaDxB8OveV1wJ+p88pE7DDazg1
VGiNRnAph0kXy5GQnRwiTkajZYvxxlXbo+FLeiS3QGqiIRr7ZkYNyO0KvnAnX56d4S6cxrEi0eym
D9dDcug9z4gykGPxOlEHH7KFJaVqePBbbmzs8//Il2u4bAaivXLzui0QqOZZ9m2ClCiVM8atXZ8N
MHsE9QzVc6XF9h3UXhNHgVfGJTYRYKv9lQCEGw9VbW2nYgpxSpxdGshAYxG0TmiTDlcJuz9jNQmk
KJi3EX8xgM7vJu5dvbOT8MYLkmvS85fscHI/bv3LPyH0txp0c329ORZ13LKZ0X+pYQ0ZM/PIU/Mx
HVGuJyyEtDsNC0Upc5JetOVlA1Jiaoj6LMlVrsxxwkS6YHeC5Fxg6BCwbkiBcn0G7RAgqJaCLDZv
wMYDFq4IOZDHxKapxULax4LlCG5Gd+0kRvy7eyqU8i1euDodam4bitWaGk88b3pUPER7qbM6IYEz
e922Y7H9m7K7O3insBY1jURFNKv/NwseqORWjeh8z3alYlyPALIEas3NZ8XaKlJZiU0az96HxTfc
SUZv/99O12m5ozR6WtIxw2TTGH3nedJOoyz6+JfMvvgq4DlQOmCVr5AgRC9QiGgZlVHPDuD5f44e
OpxelhSFg2heKuXzgV5TaO+yzMirJA7B0JjfK0/5ClBtMsl3N69TLlFjW4vNbeRg01j/0MZ/ZHNN
9ajJXdrkuFAcEuhhBFMo76HatjDDeC8WpXBnmBVNTRup6MouktUDdtNWXK7iJd6Vsm2oPrxdcp+y
pCUQ+jtJcmuJKxfsanKpwB4iy1n/8NVNmUJhi2/L5gv9ZX8Rk+BHnLSVKaa1uyRjTbqUbcpxfJSN
1xTe88Dkj/E6E60IQVwXlS6xUqshUawEQwTEFHi4xoR8+ZFQRbx6iY4ClodyoXaSOL2nlzlFXssl
xWzX2InfweQ3YhhxmoE+he9Rzy7v5U3xoRsWpz5Pa/0Hrhker87wrKl2FmqioO5ePg8lBh/aDg0E
9GG+L+blj7RZ0rfezOHlwXSQA4xqEetqDUvS8hk00dnmPqrWjGkqpbvvGUWpB3W13GANGtXgFCJz
cLzdg7bN6BWHGRkiCUUjiOaDzMwdDCrNuDt7gboLYnJif32X19IEI/D45cHgBADjcugcQcA0n/eC
p973J2ZyTl9PkXGy9kx74SMRM4B2ZsnlYo7ZXiSIbWxiYIxTpdZGfMUHIKN067HiMQTSKXs9UCf1
WtvEo0cq2HIjIpcuSXEPCt83rEi1j3aBM1nj4tDyWqxnIXtO0sa7OsxFALwIC8/hTkcexazRgG7l
BhcyXhIOA1zaUayB6NbgGw70xMgHe8lt/5Axww2JQ+csV1TccSWontBm2/NSQPQ+RnLVHMjIZBHm
y/5sTU8ZKmodwJsfgGxSo8bh5L8w8LyRjc7K8g5pjFpNYV31MYj2B9On4XJB1C9r1dHu0JbhX7fq
4buQRLh4K20PcAy5Ew6Fv1jqnUS8oM/owyEPC5KME1A5spv2GPJEbiXgv6MRjbaErR0kIEiPH/Th
fGm17GCstRtKaJhfIdZLXzqLgny4w/U89SRo8UuyD85J+3h1vrar+T27PAMi7kWgFIkdVKYIVmWt
D5zm30Mo2YJBpd9Dbg3kXD2shNOv5zKchXAr4Re5KMvTp41oi1qxifPW4xhbKjhbLnguoBDOi7Wh
R+ob380jQnYKjtRg9Gykv6ngMCBSSOm41slg3jnoKWVgOP1LeIgtsIlzA6UiFujFkw7LlTEvQ8KS
mr9pwUqYsaLAtSF5Q+gtAqzhpM5rwFH6S5luwmZ2oiifk6MjYVYEhzKZRkKjZE3jbPVKX6hnzsgM
iwRqJ0yU0b03J8IfNaGzeqQsnFcVQD8tucygNEvpO3agXPBDt8M0mL7myYdFTpephwVZ7+QHQyEZ
uTt5MnBZXK0jtoT7LDvw+t6JXvcSAP1yBSs303IMk0SMjq2gokhY9BmXyOUqBPfgPwhIjqjXUfWN
DKHK4jgZCjBIxk00KMrawmMKQhFeRWOUST92+2hrREPDxl8C3QqCRHEsfS/jFFfcwbhejm/Rcvn5
g9Q28Z2N/L/s9wU5wCLAALRsOxgGBAxMf+pFHB94iOmWT2vk3lb8IkGVvQIJzuEQtasp4Ygf0vL9
5cNu3OM80JYrTXKa5yP6yocaszKCRaEoVFSNO+2iUqkMMBpQs8Gbcd+SKACoT3dh0SLYBmOAXohj
Q+AbxEyLaqRZOtwJbED8nPjLW2pv4mm6VMb1JzvP81ZOM+cxs6STaWXo2dO0oXwPStqSjVOUfz93
f/dLAAzEgm+imVhstuKAgserF7KgooYxJwA8UAybw+usPa5LdOj2ZFfo9Er8AZopJFBvy+pqff1a
CnMUAeD5yEFVH3wyUyQKJmmEejlXkH/zuHULN63E3zA4qqqqgjtdPPZc0nIFRhDGG6SGWShnizuQ
wK7UmYHISPqS9jCj8eFIosxVCHEzAoUGD8auwPCFf5diMVhyv4dIt7o1VeiedtI2uVkZhQqZGMU5
XPbJt1EKa/1RxWSNHdW31eE19cz7ncrz7VAxBGHvOvV1Qf5yC0SiwuXfK1ibSWwd2vt2fE0ZYZVX
utnBMCaTUHx6ViKKZquvg0Xml9nKBmhR6rrvBXLRYHyi8vK0z0uzI/whTOTPV2kZLnEHclzzOTFj
OlNQQ+mvizhH2EY86B0/cBCTAYsQ/EptKu1gU8BGpEE4ymRU8xm3qgO2gfD0H24A5UPdL2iNzNaf
GLmBYAEbwyEasCAxEyIEfTg2MGh0CdDHKa11P0o65yaCf7yiu4oQ5qaSj/WMhax1uuFotBcAU2kn
Snow27gqWr6n84EkD5VsyE19HgkdHO0+T5KeNbheVwywju52eh87zTguXBhuv835F+GO7RSQQfOd
SG3UVJVLhCo/heW4X2CZmbTS7mxnPRguumiQguhytJzbHOiHpNj2cEmWEMNsymPXVEp99pUEN3zS
5mzPQ9utFl7YdhHMHMoEn4cIVi2GaSV8yx/a+Qy2mh8gblcELrPV8vZWGKDRa1t9+pKjZq8FNKC0
BStw58zaLO1CmtNQSKx4U+4CN8SzRYl+LJuyGfittEvpRsV+cCj0sTY59VzLE32sT3spYbclXA0I
uPVnPTPcn6556VcI45Hgc6JeKHpzZQOidrYtEVBaytl36uZmV9BGC5t8fpbDceOU1wlT1lZqqUk3
GSrgmHdKLhIRCAktfKsCzvvGKNQ6CGRirwcOVJCq4l/MnYXLccggr9/CyTXG+JsfkRmvawdkhWQn
5fapdxBXKelztZu6++rrtJsfTuhrISexm35dWOCiSP+ix/e0GLJEGSCyUkGS5TkuAdrQq4YuXWFQ
Ry6oaQJr4QpijXiZwL4fVI77ZTEJ+Q/LZgV2v0aeqI0QUNWfeqfPN8rZjxnt5uxukz+SDkVHoU0u
Qj5kJAtkkOmj5Xww8Svv+xHPkIq1wIVQ5XOScriwLPBGQfXvEoQ4Tkq3t2ZIkblzIxvat9+urJh8
t5kkiH1yxpZQYEzcBLHV/YQ15My4cL8//lAjVSs9rFAspyrNbKWvTSblD+qYD9GqDmbem6dDXGgo
9gl7AOoEmxV0Vw8jW6oJqB7AYez/4ouiZYEbSYQ4i1e4gujTkLmHVYCAI5ddedhlUDd9CA4bny9o
OcZnFF90Ed5Te8nWym8eNEhCKSK5AX6wt95ElwBuPA4AUFEQGweM7L1omrpDpZikz/EVUaJH9+bP
gFqezShMeh+NdlLQnB1694Tv00zSYfBpLotZS7qqH0iNNnzaz2jfwltAQoTCeM5YUBu0092ZzquD
92W0Q44vcWTMR+Co7gzReomK+NRedoQcHguqrTUYEhuDLP27674doLQeyHkUTvFneUxymkNeNKVK
kcRZwVHJ685hZDV6ccS/weWrWwglmlsCBFWV76cWZcMYL6FpB+3G1sXjVz8OqrxUith9EejFWxIX
Zdk5EbDGKRA8ZUdAJGBfnDb9lDXklfZOhoi3Tib9TQI4peb7hvix16J8yu/2due3DZNJeJ1/9/AD
uuTel11mfyC/njkAt5rqPbRSnCraT/2ExfjbHK/O0ptdobR+ZFkW6XpvJdQo9ZuX9aBj5tsVAYkl
V5UglL07ORYUVQCkzYRcASetw37ojaBxmnPqrQOUbPjEwN5pKPCpjJudQaz/Py8TdQZdaTUJy8AK
p2uiY6TyJ3N8/WvNq9IBQiHL3ekmKgb0wPYU+FoMDxNVXZgRSUaOCndee4hYePfapQaqjPsPvBsw
OIRBnOb2RAYQ2WjeY7lH24V4iOn9ixCspzCrnylnodL6fru11Y+83K3n24jBJllMDkl/zDtFm4/j
/bFTh9Tet8c7dsPebCpoTofRKopje4PF6b4N0n9ZBa3+SPQLYTN5MBWq+c/q1tYRhvuOkPniYz2j
+UCzdccWuC3JkFDhEST3Q9FCUl+8AAoUTtU+awSuQZT2XVB/yvBInVS9IJteheUW7jM3vYfVTJWZ
iJVeHbbty41RqaAdYRW9G3B91JSNHhgk9lVyFlG7L8FKYSLf2o7OiWKnglfaQZwtsj0CzdeYxbgB
Dwg9w09kNMN3l3J2Rd8QKvS4Zrf7nP2/u5PmGKhre0mY5ClyRcBpXBxAPT6k8S3GPOYNgOaGCT5j
9HAi/mDMVWaA2FFjf7qCxMpETHtXMI0LdTIe/sbJ/8AoL0wVPs/5SVnD2giIPpM71vVLetcTqSv4
FrofuvPgc6OEiwUv10as0H57wD/Cg6koxqxCXYIaaizjFgBcAPYqEitwRJCvJOfTswPM3huF7AWU
ZY2A9gI2fn8ZCV8+pv6GS5n7ndfduCR4lqbW0WvtzKUGQzwmu20mYecsNNdIz0CKYuvjB3NqpYnm
uUkJPIrTjeq+u3CoCIp3IVX1CjGdfvalcHA6hCEJy8dTzyJ1v3IKG0bmhjY8CfdzGWd3BLw4q+uV
Pnr9QKNXZI8SwA44uOtilw0yubO8reCzynqICwf01CQCoOBAgjau/EtXxEa4cHIDgcUK9afvh2gN
rR0q6zJ1CvHgH3ii6Khi0Vd5aimejnv7nhZDiwh3CjL5YERzKVR7UXXfYpTsMtIv9sN+KTP53Zbu
Qkk2PfX7dEXZKzhT8sYGxERExkZkcQvcwmpasZdk2VP7BMqAiZ47acr3vuEcKMWuOxyw78yp7JPE
7+sYLxb1u7NsgdxU5FEW3M47uLx8nCr+grQxs77DylzxQvvxJ/261+E2iU5M2eqZPzWn8EjASSsP
sTJhQ3lfHvC4OrTDj331fk0up6o2qcMuBWZ1ECEp/7YVzWg5s/qNty+fa9mSalGIVwwxKNlFbKaZ
v8fB0GC391vt2Z9x8U73P7Xcd0EAdfUW9c1o1jpJssj++0tHsSh+xlJb+fJATRz6H1FdbsUK+/Jf
xHiqx9UHXOMxP2cCQ6+2uW+vdDJwdn4HQjteC/lP4Bkm93NQzbwl1w24ylRPF2Vv6UmsGqTKJHAR
5DGeOeT8APTBK67oRNd+l3ZmP/9Z34BltEksrDGd0KDJm/oFulYh6ELRaSs6RxbI+dwfg4hu7qxm
/QIu95Rk0AjsJ6EdmcneJAICmZ77S3AHtYUSw5X+j6jmsgONB8pGeyVVhIG0KfjzLZq24gaheqXz
wK1cytm4tYFcM1nsm5KRxxlvk2o7drPlFzf0WBGPmjeccxZWBIQ9piy2TsCGH7og0hNOimx0EGsI
i7DFvHa7v9taXVO+8LizuqTjjb/bCYoJGb+kTpZHSl2nngkh9vHJ0mfKpo8m1zAKX0eT9KeqTq7H
B1/0zZtUuhe21p+qT1LO/5XqKxpmWEwskPWhI3TjAhrA/VPveZjtEp+iSJ7uUiiOowOqIc6OMbSP
RK8kMbngRD98IdR61ruwy7ATXf6rN19Jw/jGakkX+GwAPtpv+5r/tm/AXQBljAzl2tLz432oURVh
yqfmiPXrzrrGa4+gwclI6fNGdxEAR61Y+54Mip6C3FLMHD+9jErTwlwq1vjid9sysOuArfJwKkHU
g3rVJQXuFljE1Ok6nFk/toaMeq9oKnBK1B9bhOJn65MhNw+Bio/Daz0Nm/PKycg95Z27wJ0t0ieA
cNtGyTrFpu/AWw4ZhpX/jRj0gGMrF5dWObt8MPeeGmtgOma20tRazK9lNCPLU7vriMHZC9Y9YYoU
uEqyfrY0o0HlTw3fiU/0zTdt5DXCY2tyiFXKPRk0W/N2YolUZlOkIyoniIy7ulolpnJZ4CNhdQoP
tcBICjQMYxRePUSs4j54D3XHRw58R6bY725ITtp9+s1YtOTTrafEZbnhYjDJLoHHeeVhbEOqMnpk
4tewseA9d+qC7pQqueWILWVBuY4ReQh8SmSPNtFAzR3DHy8z/vjRvv0JVPLe10z5rVR1TYqPddFD
Fkwrqv1U2l6qUkMC07dLV1CY+DaFm/wU7TVzoWP87ZWt6upk3AbkpKXDQolsXNy80idO9MLOVPUa
cgthpZNDgZ9IN9RQ0uxsIXFZ21o6IjmuNXe35iwcn8rd6kmMsx95dex51qlBurKQNZ5BSGrZo+mu
ykkfCA/kZlB6/0hUjLj6kaZTAshGyjsgnDB2C9iMqKQzSqcIynvMs5uWyr+32F/AvKQzaSgZI9C4
PSNSmGoikZtK6naUfV7uB5X4ev/l1VxVM6f64PGrHeAz7etZWqRWR3SF45tAnVQHc1fQpY61xI7Z
sqmzjx4EUtnGvXcQ24aRgikRqcCxRkZegdRa/IBfuUzuwxJgtJGKw1XIWLCpCnOZ/KiEppPabkEw
XBijoBWnUiF69H1UcqRzS5DdN733u/y/zNhisDGZLRXYUk9xhFUUklgOn0oQ/Il5IR1/DSDTCjEc
UiEEDI5aJ7GjSIDCYE4zBFKx+Lno+9t697VofEMIB9xqRwS9Xoj9gDEUeD5VyYenVi3lEO0/rXyD
KF5fhaN/jzgHoYRyQH06ewjD7fKnLFR+zMCMkvWJ3X5BkLXSksMPhpErcmiC/MKs+UsQQuNnGqMb
dXeehq8am1Y0mqH+L++g3XiLjBRKtxMYbgYT0+OW5Kc5aJOIBHAW2SLcIS5xa/bcxb6YJ0ggkeKV
LgrwP55OW/jhEk98BeTwrd10DdQN+byeYDMiMhynVmxc2IvOlRVch33rJ0qYRedoKNwX88c8PXl8
ss9vyeUfq+ACYQTtGiNOaVNw6z+pZTjgf5odAmVw/GhStPJpmz8/0P8vbGT8vVLszD6xSLBp2UQM
xIcC+kyfIQ6ymyVWEFtPoDCBoVz1haOTW9y1jSEeBnxIJcmgCEWUjrU48+2l0y2jYlwdsw/WUZGy
rq71m8mwmCkFFPK6nCTCOqMeoKM/wgxeJfruc8IO2OZQ5HXZNyWYZXr2/DIiv5GyEhUDGGNOA6gS
aBi7k8mESwTJMB2V7+u7cKCB3MRTh7rNehKLr5Jy8i3aSiuku31E3u7GDBIjptJphk/ZSP+bCR2T
rN7GPF6OyclV+2AKMsQaaeq4De3y9VrsT7UYQQ5m3nH7G2IBWp3vJOGSb4WGHP3e9DKzrTZU2bIq
mw99K2A2ce6cmgwfacIT5QJAWpxo2n3ShynqKZGGtBleRKe3FjF3ZkSDazxN/a6ncK2YZjrAp4U+
WN0Dcwhr1XBhvxpEC9aQ5ZD4usX8tNZs2dRZfiV3EXGrdkC5Mrh1QatgLYvLS+/ZLCR1NfyRtAO0
qNAX1VHSakalLwyN5L7HbdnMbM+WNTLoih0/WYWRWx3GSBo9YUUzAggNJ7F1a2/XMf+w8bCP2vEF
uZhrLaBXRl+0bfMdav8WhBlGYVJbEgs8y2AnMOtii7DvOcvZRmcOjgLO9pji1LWM1yUfkFRWV1kb
m/TzUDUzOuDJo4Be5bvCFf9fPiJ48s98gbOujvfaagKuyuYZaHu7auonhuTfVv5ohdu/3upo6hZy
kGOg1bVVeNVNshIWBM5wRb5Z1eFApHi0RCljmXSG4egz0vokrv5wCPC1cYDab0x0r/cDpeGhHL7P
565p6xpAsWzBaOKAQLakmuwtXd7jc7tChOqYyZhQt/LUUMrN1U2AuBWFfaiG+lFvqWw4d59gwMd4
27d1svvkzI36T2dqPG6z8VP7iS7Bq+4OZUfJggT9UJjDdSSCvrJrx1N+U9tLZP7IdVlMdiUyge9d
hlIFfyw7lcgyJg4iHpajE4rrcDtWs7rhe6xhH8bZVmif17XQnBq+eCWdQT1c3JKW9VCwKobc5j2y
O2T3hSmCnCrWNuVNrDeIrNl0QO/ADC4ogDOVFFQFlo2gq4DSocn6gnkr0VI2b2m30f+hQ+IdQrGn
vjakqzOy7DeEWjOeJNzb3rE90MKWSWHFHIGfvSuA7BxSw5AcxS4AxtmJG3zAOGQhUm3AGI070Zhu
2osWz+r/dOQVQWknTCkgusFfWlWvS/1yKS45Iau4UcN9IoKe/XTI8AZnzTG5ijseyNmrjrydJVhd
7adKj1uCmquz/w47wBqwzekuLCx3D5OB7glvtfc0TybfH4UTTmzVsBcRx+hRqoN+hViMxPCXh6f0
yUZS+eUtVOAut4/1Mp1zOrsIVTVg+yaxmMuhyzIG8qpyJcrraAumGjyFNm1ntQE353Gwgk7cARr6
j2apdnYcG2obX+rYPVUgUqwpvUhFyGHzMp6mS+ZmEl/wdNYYy64oFYozqWJr4/LOCwxZAHpNvCpR
7niSPBZRejCQMSzJyN2aTo6UxCr+urVsuTj722mO3xV1q65uGp12F7/uFRKSLEBT41LvdVy7i5Oz
BfyAmnZ29yw5uvLGFVWkklG/HxzeIeRryIqlUlLsZZ0GnLJluj6sWdZWFvBnt8ZPTncAkBALURU7
XGHE72BrnZPS4Bbz9itcZaOx+4L30Z5rCE1RuDZi98cmapgD0x2GQTgo/Mespa2BIoqrUQnhBaDB
RSXIIfD/lSQwlmMXaAo73fAUHHAIeREaHEHOAiqRXnLlFQMR3SRqoF9x8OknLqUU3S/huMiSZDpn
OX0t7PseBEMcuCTr1mpEc2xfcIbaBp39t8maF367SWPGMDBypk5rWPPU5DB7mYxwnAmCRHGBigH3
OuuHT0UkzsRXJQCCWuizgrcLc/FpzHy3gd20pxreFWPoXjI2XTn29k4ziFXvOmRlVe5Vllmn7VEo
5rC331JBqDrlogBvTS0cEJtYVEjKoKfFHk+/2heGCJx65UCTFvOPvJn+svoXRewPGPu8PLF0tXSH
lzBI9VoN3tnbSHYy0lOjoiK6AJpRZP/0bHkDkgHs2GxwM3hvb45CUdG9P1G017BbTIb7tAL2R1t6
8VoGfZn4vJJvjLFFfmfWnRiiv5J2NZGZtjGhaYI6+DDxqirO8AleQC3bTTPlnWrYG42ZioMfkE35
nmqlk6mT8/4CUQYvtxJoDcohycNJPOR8T+JpotTsGgbnJ78Y+ow4PRayJYnxGMrwRwBMtTVsE2ax
xpFLh2EzYg4rDsE7bYYB04WnpVoNwIV+SPpliEGPnZn0i6KV/rGkHTYWIpb8XN4jvpLtB9g4bp/6
lQXNHvwYfLwJv+Sy9NBEQII/P3jO986/UzxeN+ELF1mSL2aecyBslcDgCqR5mCEWkwnh6/q42bxj
cV2sGMXkItDJ2Pk+/+fEATUUiwmmpj9kHgziYL7PNbhH8tx2UxKRsU4EbX0rLVFQ6vVAFtScaTUs
CkyroHHnVQ4CND8/KiWX0ABfwZLELoYEAeF8VeZ3Ixq01Z+iieYzHpCE4rmljtnKo2QsxWBemOG7
PV8s/9YvLTuwT4+P5OvidBvZMlcxlaf53bv7CrLdHvWH2mtLNTB15bXIARHz1gXQV2RufGsR2mP7
cbhHPNju0q7LjNWNkIk+yr08mam52Wxof7s/avdCZQTLfwZJ5JoMhNfB/Jh4ZQZrJFcXIQ1vzMiD
PlNUR0LbGLST0OsJKDqJ/P/BSXsTUFKrozA4A33xqueDCzSB57Q3tfuveW1M9uE/3ym1WHWe0Ksh
6Z29H44p9ZLyEwMtv1i3xt9/ENBXf423uiTEsxrfgcSi6rA0wZwmXvfE5TuOCgBauT43SDa0ZGid
4fb/H9j7EqE=
`protect end_protected
