`define DEBUG

module eth_encap #(
	parameter KEY_SIZE = 96,
	parameter VAL_SIZE = 32
)(
	input  wire        clk156,
	input  wire        eth_rst,
	output wire [ 7:0] debug,

	output wire [KEY_SIZE-1:0] in_key,
	output wire [3:0]          in_flag,
	output wire                in_valid,
	input  wire                out_valid,
	input  wire [3:0]          out_flag,

	input  wire        s_axis_rx0_tvalid,
	input  wire [63:0] s_axis_rx0_tdata,
	input  wire [ 7:0] s_axis_rx0_tkeep,
	input  wire        s_axis_rx0_tlast,
	input  wire        s_axis_rx0_tuser,

	input  wire        m_axis_tx0_tready,
	output wire        m_axis_tx0_tvalid,
	output wire [63:0] m_axis_tx0_tdata,
	output wire [ 7:0] m_axis_tx0_tkeep,
	output wire        m_axis_tx0_tlast,
	output wire        m_axis_tx0_tuser,

	input  wire        s_axis_rx1_tvalid,
	input  wire [63:0] s_axis_rx1_tdata,
	input  wire [ 7:0] s_axis_rx1_tkeep,
	input  wire        s_axis_rx1_tlast,
	input  wire        s_axis_rx1_tuser,

	input  wire        m_axis_tx1_tready,
	output wire        m_axis_tx1_tvalid,
	output wire [63:0] m_axis_tx1_tdata,
	output wire [ 7:0] m_axis_tx1_tkeep,
	output wire        m_axis_tx1_tlast,
	output wire        m_axis_tx1_tuser
);

localparam TX_IDLE = 2'b00,
           TX_HDR  = 2'b01,
           TX_DATA = 2'b10,
           TX_WAIT = 2'b11;

reg [15:0] tx_count, tx_count_next;
reg [ 1:0] tx_state, tx_state_next;
reg [15:0] wait_cnt, wait_cnt_next;

//always @ (posedge clk156) begin
//	if (eth_rst) begin
//		tx_state <= TX_IDLE;
//		tx_count <= 0;
//		wait_cnt <= 0;
//	end else begin
//		tx_state <= tx_state_next;
//		tx_count <= tx_count_next;
//		wait_cnt <= wait_cnt_next;
//	end
//end
//
//always @ (*) begin
//	tx_state_next = tx_state;
//	tx_count_next = tx_count;
//	wait_cnt_next = wait_cnt;
//
//	case(tx_state)
//		TX_IDLE: begin
//			if (m_axis_tready) begin
//				tx_state_next = TX_HDR;
//				tx_count_next = 0;
//			end
//		end
//		TX_HDR: begin
//			if (m_axis_tready) begin
//				tx_count_next = tx_count + 1;
//				if (tx_count == 9) begin
//					tx_state_next = TX_WAIT;
//				end
//			end
//		end
//		TX_DATA: begin
//			if (m_axis_tready && m_axis_tlast) begin
//				tx_state_next = TX_WAIT;
//			end else if (m_axis_tready) begin
//				tx_count_next = tx_count + 1;
//			end
//		end
//		TX_WAIT: begin
//			wait_cnt_next = wait_cnt + 1;
//			if (wait_cnt == 16'hffff) begin
//				tx_state_next = TX_IDLE;
//				wait_cnt_next = 16'h0000;
//			end
//		end
//		default: tx_state_next = TX_IDLE;
//	endcase
//end
//
//assign m_axis_tkeep = (tx_state == TX_HDR) ? 8'b1111_1111 : 8'b0000_0000;

//always @ (*) begin
//	if (tx_state == TX_HDR) begin
//		case (tx_count)
//			default: m_axis_tkeep = 8'b1111_1111;
//		endcase
//	end else if (tx_state == TX_DATA) begin
//		m_axis_tkeep = 8'b1111_1111;//dout[73:66];
//	end
//end

//always @ (*) begin
//	m_axis_tdata = 64'd0;
//	if (tx_state == TX_HDR) begin
//		case (tx_count)
//			16'h0: m_axis_tdata = 64'h11_00_d1_91_5d_ba_e2_90;
//			16'h1: m_axis_tdata = 64'h00_45_00_08_55_44_33_22;
//			16'h2: m_axis_tdata = 64'h11_40_00_00_00_00_2e_00;
//			16'h3: m_axis_tdata = 64'ha8_c0_01_64_a8_c0_62_31;
//			16'h4: m_axis_tdata = 64'h1a_00_76_37_76_37_0b_64;
//			16'h5: m_axis_tdata = 64'h3d_00_00_00_00_20_00_00;
//			16'h6: m_axis_tdata = 64'hFF_FF_FF_FF_FF_FF_FF_FF;
//			16'h7: m_axis_tdata = 64'h00_40_00_C0_00_00_00_00;
//			16'h8: m_axis_tdata = 64'h01_08_00_00_00_00_70_00;
//			16'h9: m_axis_tdata = 64'haa_aa_aa_aa_00_00_00_00;
//			default: m_axis_tdata = 64'h22222222_00000000;
//		endcase
//	end 
//end
//
//assign m_axis_tlast  = (tx_state == TX_HDR && tx_count == 9);
//assign m_axis_tuser  = 1'b0;
//assign m_axis_tvalid = (tx_state == TX_HDR || tx_state == TX_DATA);

/*
 *  RX path
 */
localparam ETH_FTYPE_IP  = 16'h0800;
localparam IP_PROTO_UDP  = 8'h11,
           IP_PROTO_ICMP = 8'h01;
localparam ICMP_PORT_UNREACH = 8'h03;
localparam ICMP_DEST_UNREACH = 8'h03;
localparam DNS_SERV_PORT__   = 16'd53;
localparam DEBUG_SERV_PORT__ = 16'd12345;
`ifdef DEBUG
localparam DNS_SERV_PORT = DEBUG_SERV_PORT__;
`else
localparam DNS_SERV_PORT = DNS_SERV_PORT__;
`endif /* DEBUG */
localparam DNS_PARAM_RESPONSE = 1'b1,
           DNS_PARAM_REQUEST  = 1'b0;

localparam STATUS_SUSPECT = 2'b01,
           STATUS_ARREST  = 2'b10,
           STATUS_FILTERE = 2'b11;


/* general regs for parsering */
reg  [9:0] rx_cnt0, rx_cnt1;
reg  [7:0] hit_cnt;
/* regs for parsering */
reg [15:0] rx0_ftype;
reg  [7:0] rx0_ip_proto;
reg [15:0] rx0_dst_uport, rx0_src_uport;
reg [31:0] rx0_dst_ip,    rx0_src_ip;
reg  [7:0] rx0_icmp_type, rx0_icmp_code;
reg [15:0] rx1_ftype;
reg  [7:0] rx1_ip_proto;
reg [15:0] rx1_dst_uport, rx1_src_uport;
reg [31:0] rx1_dst_ip,    rx1_src_ip;
reg  [7:0] rx1_icmp_type, rx1_icmp_code;
reg [ 7:0] filter_ip_proto;
reg [31:0] filter_src_ip, filter_dst_ip;
reg [15:0] filter_dst_udp, filter_len_udp, filter_qid_dns, filter_src_udp;
reg [15:0] filter_parm_dns, filter_qcnt_dns, filter_acnt_dns, filter_auth_dns;
reg [15:0] suspect_parm_dns, suspect_qcnt_dns, suspect_acnt_dns,suspect_auth_dns;
reg [15:0] suspect_qid_dns;
reg  [7:0] filter_iph_len;
reg [15:0] filter_ipd_len;
/* DB Request Registers */
reg [3:0] db_op0, db_op1;
/* pipelined stages */
reg  [1+1+8+64-1:0] pipe_stg0_0, pipe_stg0_1, pipe_stg0_2, pipe_stg0_3;
reg  [1+1+8+64-1:0] pipe_stg0_4, pipe_stg0_5, pipe_stg0_6, pipe_stg0_7;
wire [1+1+8+64-1:0] pipe_in_stage0 = {s_axis_rx0_tvalid, s_axis_rx0_tdata, 
						s_axis_rx0_tkeep, s_axis_rx0_tlast}; 
wire        p0_axis_tvalid, p0_axis_tlast;
wire [ 7:0] p0_axis_tkeep;
wire [63:0] p0_axis_tdata;
assign {p0_axis_tvalid, p0_axis_tdata, p0_axis_tkeep, p0_axis_tlast} = pipe_stg0_7;

reg  [1+1+8+64-1:0] pipe_stg1_0, pipe_stg1_1, pipe_stg1_2, pipe_stg1_3;
reg  [1+1+8+64-1:0] pipe_stg1_4, pipe_stg1_5, pipe_stg1_6, pipe_stg1_7;
wire [1+1+8+64-1:0] pipe_in_stage1 = {s_axis_rx1_tvalid, s_axis_rx1_tdata, 
						s_axis_rx1_tkeep, s_axis_rx1_tlast}; 
wire        p1_axis_tvalid, p1_axis_tlast;
wire [ 7:0] p1_axis_tkeep;
wire [63:0] p1_axis_tdata;
assign {p1_axis_tvalid, p1_axis_tdata, p1_axis_tkeep, p1_axis_tlast} = pipe_stg1_7;
wire filter_mode  = rx1_ftype     == ETH_FTYPE_IP      && 
                    rx1_ip_proto  == IP_PROTO_ICMP     &&
                    rx1_icmp_type == ICMP_DEST_UNREACH &&
                    rx1_icmp_code == ICMP_PORT_UNREACH;
wire suspect_mode = rx0_ftype     == ETH_FTYPE_IP      &&
                    rx0_ip_proto  == IP_PROTO_UDP      &&
                    rx0_src_uport == DNS_SERV_PORT;
reg  filtered;
wire filter_block = filtered || (out_valid && out_flag[2:1] == 2'b10);

always @ (posedge clk156) begin
	if (eth_rst) begin
		rx_cnt0          <= 0;
		rx_cnt1          <= 0;
		hit_cnt          <= 0;
		rx0_ip_proto     <= 0;
		rx0_src_ip       <= 0;
		rx0_dst_ip       <= 0;
		rx0_src_uport    <= 0;
		rx0_dst_uport    <= 0;
		rx0_ftype        <= 0;
		rx0_icmp_type    <= 0;
		rx0_icmp_code    <= 0;
		rx1_ip_proto     <= 0;
		rx1_src_ip       <= 0;
		rx1_dst_ip       <= 0;
		rx1_src_uport    <= 0;
		rx1_dst_uport    <= 0;
		rx1_ftype        <= 0;
		rx1_icmp_type    <= 0;
		rx1_icmp_code    <= 0;
		filter_ip_proto  <= 0;
		filter_src_ip    <= 0; 
		filter_dst_ip    <= 0; 
		filter_dst_udp   <= 0; 
		filter_len_udp   <= 0; 
		filter_qid_dns   <= 0; 
		filter_src_udp   <= 0;
		filter_parm_dns  <= 0; 
		filter_qcnt_dns  <= 0; 
		filter_acnt_dns  <= 0; 
		filter_auth_dns  <= 0;
		suspect_qid_dns  <= 0; 
		suspect_parm_dns <= 0; 
		suspect_qcnt_dns <= 0; 
		suspect_acnt_dns <= 0; 
		suspect_auth_dns <= 0;
		db_op0           <= 0;
		db_op1           <= 0;
		filtered         <= 0;
		pipe_stg0_0      <= 0;
		pipe_stg0_1      <= 0;
		pipe_stg0_2      <= 0;
		pipe_stg0_3      <= 0;
		pipe_stg0_4      <= 0;
		pipe_stg0_5      <= 0;
		pipe_stg0_6      <= 0;
		pipe_stg0_7      <= 0;
		pipe_stg1_0      <= 0;
		pipe_stg1_1      <= 0;
		pipe_stg1_2      <= 0;
		pipe_stg1_3      <= 0;
		pipe_stg1_4      <= 0;
		pipe_stg1_5      <= 0;
		pipe_stg1_6      <= 0;
		pipe_stg1_7      <= 0;
	end else begin
		/* Pipelining  */
		pipe_stg0_0 <= pipe_in_stage0;
		pipe_stg1_0 <= pipe_in_stage1;
		if (!filter_block) begin
			pipe_stg0_1 <= pipe_stg0_0;
			pipe_stg0_2 <= pipe_stg0_1;
			pipe_stg0_3 <= pipe_stg0_2;
			pipe_stg0_4 <= pipe_stg0_3;
			pipe_stg0_5 <= pipe_stg0_4;
			pipe_stg0_6 <= pipe_stg0_5;
			pipe_stg0_7 <= pipe_stg0_6;
			pipe_stg1_1 <= pipe_stg1_0;
			pipe_stg1_2 <= pipe_stg1_1;
			pipe_stg1_3 <= pipe_stg1_2;
			pipe_stg1_4 <= pipe_stg1_3;
			pipe_stg1_5 <= pipe_stg1_4;
			pipe_stg1_6 <= pipe_stg1_5;
			pipe_stg1_7 <= pipe_stg1_6;
		end else begin // Zero is inserted in regs.
			pipe_stg0_1 <= 0;
			pipe_stg0_2 <= 0;
			pipe_stg0_3 <= 0;
			pipe_stg0_4 <= 0;
			pipe_stg0_5 <= 0;
			pipe_stg0_6 <= 0;
			pipe_stg0_7 <= 0;
			pipe_stg1_0 <= 0;
			pipe_stg1_1 <= 0;
			pipe_stg1_2 <= 0;
			pipe_stg1_3 <= 0;
			pipe_stg1_4 <= 0;
			pipe_stg1_5 <= 0;
			pipe_stg1_6 <= 0;
			pipe_stg1_7 <= 0;
		end

		/* DB reply */
		if (out_valid && out_flag[2:1] == 2'b10)
			filtered <= 1;

		/* Packet Parser */
		if (s_axis_rx0_tvalid) begin
			if (s_axis_rx0_tlast)
				rx_cnt0 <= 0;
			else
				rx_cnt0 <= rx_cnt0 + 1;
			case (rx_cnt0)
				0: begin // Reset all registers
					rx0_ip_proto      <= 0;
					rx0_src_ip        <= 0;
					rx0_dst_ip        <= 0;
					rx0_src_uport     <= 0;
					rx0_dst_uport     <= 0;
					rx0_ftype         <= 0;
					rx0_icmp_type     <= 0;
					rx0_icmp_code     <= 0;
					suspect_qid_dns  <= 0; 
					suspect_parm_dns <= 0; 
					suspect_qcnt_dns <= 0; 
					suspect_acnt_dns <= 0; 
					suspect_auth_dns <= 0;
					db_op0           <= 0;
					filtered         <= 0;
				end
				1: rx0_ftype <= {s_axis_rx0_tdata[39:32], s_axis_rx0_tdata[47:40]};
				2: rx0_ip_proto <= s_axis_rx0_tdata[63:56];
				3: begin
					rx0_src_ip <= {s_axis_rx0_tdata[23:16],
					              s_axis_rx0_tdata[31:24],
					              s_axis_rx0_tdata[39:32],
					              s_axis_rx0_tdata[47:40]};
					rx0_dst_ip[31:16] <= {s_axis_rx0_tdata[55:48],
					                     s_axis_rx0_tdata[63:56]};
				end
				4: begin
					rx0_dst_ip[15: 0] <= {s_axis_rx0_tdata[ 7: 0],
                                         s_axis_rx0_tdata[15: 8]};
					if (rx0_ftype == ETH_FTYPE_IP && 
							rx0_ip_proto == IP_PROTO_UDP) begin
							rx0_src_uport <= {s_axis_rx0_tdata[23:16], 
							                  s_axis_rx0_tdata[31:24]};
							rx0_dst_uport <= {s_axis_rx0_tdata[39:32], 
							                 s_axis_rx0_tdata[47:40]};
					end
				end
				5: if (suspect_mode) begin
					suspect_qid_dns <= {s_axis_rx0_tdata[23:16],
					                    s_axis_rx0_tdata[31:24]};
					suspect_parm_dns <= {s_axis_rx0_tdata[39:32],
                                         s_axis_rx0_tdata[47:40]};
					suspect_qcnt_dns <= {s_axis_rx0_tdata[55:48],
					                     s_axis_rx0_tdata[63:56]};
				end                          
				6: if (suspect_mode) begin
					suspect_acnt_dns <= {s_axis_rx0_tdata[ 7: 0],
					                     s_axis_rx0_tdata[15: 8]};
					suspect_auth_dns <= {s_axis_rx0_tdata[23:16],
					                     s_axis_rx0_tdata[31:24]};
				end
				default : ;
			endcase
			/* Debug Logic */
			if (rx0_ftype == ETH_FTYPE_IP && 
					rx0_ip_proto  == IP_PROTO_UDP  &&
					rx0_dst_uport == DNS_SERV_PORT &&
					s_axis_rx0_tlast)
				hit_cnt[3:0] <= hit_cnt[3:0] + 1;
			if (filter_mode)
				hit_cnt[4]  <= 1;
			if (suspect_mode)
				hit_cnt[5]  <= 1;
			if (suspect_mode && suspect_parm_dns[0] == DNS_PARAM_RESPONSE &&
				rx_cnt0 == 10'd6) begin
				db_op0 <= 4'b0011;
				hit_cnt[6] <= 1;
			end
		end
		// Port 1
		if (s_axis_rx1_tvalid) begin
			if (s_axis_rx1_tlast)
				rx_cnt1 <= 0;
			else
				rx_cnt1 <= rx_cnt1 + 1;
			case (rx_cnt1)
				0: begin // Reset all registers
					rx1_ip_proto      <= 0;
					rx1_src_ip        <= 0;
					rx1_dst_ip        <= 0;
					rx1_src_uport     <= 0;
					rx1_dst_uport     <= 0;
					rx1_ftype         <= 0;
					rx1_icmp_type     <= 0;
					rx1_icmp_code     <= 0;
					filter_ip_proto  <= 0;
					filter_src_ip    <= 0; 
					filter_dst_ip    <= 0; 
					filter_dst_udp   <= 0; 
					filter_len_udp   <= 0; 
					filter_qid_dns   <= 0; 
					filter_src_udp   <= 0;
					filter_parm_dns  <= 0; 
					filter_qcnt_dns  <= 0; 
					filter_acnt_dns  <= 0; 
					filter_auth_dns  <= 0;
					db_op1           <= 0;
					filtered         <= 0;
				end
				1: rx1_ftype <= {s_axis_rx1_tdata[39:32], s_axis_rx1_tdata[47:40]};
				2: rx1_ip_proto <= s_axis_rx1_tdata[63:56];
				3: begin
					rx1_src_ip <= {s_axis_rx1_tdata[23:16],
					              s_axis_rx1_tdata[31:24],
					              s_axis_rx1_tdata[39:32],
					              s_axis_rx1_tdata[47:40]};
					rx1_dst_ip[31:16] <= {s_axis_rx1_tdata[55:48],
					                      s_axis_rx1_tdata[63:56]};
				end
				4: begin
					rx1_dst_ip[15: 0] <= {s_axis_rx1_tdata[ 7: 0],
                                         s_axis_rx1_tdata[15: 8]};
					if (rx1_ftype == ETH_FTYPE_IP 
						&& rx1_ip_proto == IP_PROTO_ICMP) begin
							rx1_icmp_type <= s_axis_rx1_tdata[23:16];
							rx1_icmp_code <= s_axis_rx1_tdata[31:24];
					end
				end
				5: if (filter_mode) begin
					filter_iph_len <= s_axis_rx1_tdata[23:16];
					filter_ipd_len <= {s_axis_rx1_tdata[39:32],
                                       s_axis_rx1_tdata[47:40]};
				end 
				6: if (filter_mode) begin
					filter_ip_proto      <= s_axis_rx1_tdata[31:24];
					filter_src_ip[31:16] <= {s_axis_rx1_tdata[55:48],
					                         s_axis_rx1_tdata[63:56]};
				end 
				7: if (filter_mode) begin
					filter_src_ip[15:0] <= {s_axis_rx1_tdata[ 7: 0],
					                        s_axis_rx1_tdata[15: 8]};
					filter_dst_ip       <= {s_axis_rx1_tdata[23:16],
					                        s_axis_rx1_tdata[31:24],
					                        s_axis_rx1_tdata[39:32],
					                        s_axis_rx1_tdata[47:40]};
					filter_src_udp      <= {s_axis_rx1_tdata[55:48],
					                        s_axis_rx1_tdata[63:56]};
				end
				8: if (filter_mode) begin
					filter_dst_udp      <= {s_axis_rx1_tdata[ 7: 0],
					                        s_axis_rx1_tdata[15: 8]};
					filter_len_udp      <= {s_axis_rx1_tdata[23:16],
					                        s_axis_rx1_tdata[31:24]};
					filter_qid_dns      <= {s_axis_rx1_tdata[55:48],
					                        s_axis_rx1_tdata[63:56]};
				end
				9: if (filter_mode) begin
					filter_parm_dns      <= {s_axis_rx1_tdata[ 7: 0],
					                         s_axis_rx1_tdata[15: 8]};
					filter_qcnt_dns      <= {s_axis_rx1_tdata[23:16],
					                         s_axis_rx1_tdata[31:24]};
					filter_acnt_dns      <= {s_axis_rx1_tdata[39:32],
					                         s_axis_rx1_tdata[47:40]};
					filter_auth_dns      <= {s_axis_rx1_tdata[55:48],
					                         s_axis_rx1_tdata[63:56]};
				end
				default : ;
			endcase
			if (filter_mode && filter_parm_dns[0] == DNS_PARAM_RESPONSE &&
				rx_cnt1 == 10'd10) begin
				db_op1 <= 4'b0101;
				hit_cnt[7] <= 1;
			end
		end
	end
end


wire [1:0] status = suspect_mode ? db_op0[2:1] : 
                    filter_mode  ? db_op1[2:1] : 2'd0;
assign in_flag = suspect_mode ? db_op0 : 
                 filter_mode  ? db_op1 : 4'd0;
assign in_valid = (suspect_mode && rx_cnt0 == 10'd7) || 
                  (filter_mode  && rx_cnt1 == 10'd11);

//assign in_key = (status == STATUS_SUSPECT) ? {rx_src_ip, rx_dst_ip, 
//                                              rx_dst_uport , 16'd0}  :
//                (status == STATUS_ARREST)  ? {filter_src_ip, filter_dst_ip, 
//                                              filter_dst_udp, 16'd0} : 0;
assign in_key = (suspect_mode) ? {rx0_src_ip, rx0_dst_ip, 
                                  rx0_dst_uport , 16'd0}  :
                (filter_mode)  ? {filter_src_ip, filter_dst_ip, 
                                  filter_dst_udp, 16'd0} : 0;

assign debug = hit_cnt;

/*
 * Loopback FIFO for packet mode
 */
axis_data_fifo_0 u_axis_data_fifo0 (
  .s_axis_aresetn      (!eth_rst),     // input wire s_axis_aresetn
  .s_axis_aclk         (clk156),       // input wire s_axis_aclk

  .s_axis_tvalid       (p0_axis_tvalid),// input wire s_axis_tvalid
  .s_axis_tready       (),             // te s_axis_tready
  .s_axis_tdata        (p0_axis_tdata), // input wire [63 : 0] s_axis_rx0_tdata
  .s_axis_tkeep        (p0_axis_tkeep), // input wire [7 : 0] s_axis_tkeep
  .s_axis_tlast        (p0_axis_tlast), // input wire s_axis_tlast
  .s_axis_tuser        (1'b0), // input wire [0 : 0] s_axis_tuser

  .m_axis_tvalid       (m_axis_tx0_tvalid),// output wire m_axis_tvalid
  .m_axis_tready       (m_axis_tx0_tready),// input wire m_axis_tready
  .m_axis_tdata        (m_axis_tx0_tdata), // output wire [63 : 0] m_axis_tdata
  .m_axis_tkeep        (m_axis_tx0_tkeep), // output wire [7 : 0] m_axis_tkeep
  .m_axis_tlast        (m_axis_tx0_tlast), // output wire m_axis_tlast
  .m_axis_tuser        (m_axis_tx0_tuser), // output wire [0 : 0] m_axis_tuser
  .axis_data_count     (),        // output wire [31 : 0] axis_data_count
  .axis_wr_data_count  (),  // output wire [31 : 0] axis_wr_data_count
  .axis_rd_data_count  ()  // output wire [31 : 0] axis_rd_data_count
);

axis_data_fifo_0 u_axis_data_fifo1 (
  .s_axis_aresetn      (!eth_rst),     // input wire s_axis_aresetn
  .s_axis_aclk         (clk156),       // input wire s_axis_aclk

  .s_axis_tvalid       (p1_axis_tvalid),// input wire s_axis_tvalid
  .s_axis_tready       (),             // te s_axis_tready
  .s_axis_tdata        (p1_axis_tdata), // input wire [63 : 0] s_axis_rx0_tdata
  .s_axis_tkeep        (p1_axis_tkeep), // input wire [7 : 0] s_axis_tkeep
  .s_axis_tlast        (p1_axis_tlast), // input wire s_axis_tlast
  .s_axis_tuser        (1'b0), // input wire [0 : 0] s_axis_tuser

  .m_axis_tvalid       (m_axis_tx1_tvalid),// output wire m_axis_tvalid
  .m_axis_tready       (m_axis_tx1_tready),// input wire m_axis_tready
  .m_axis_tdata        (m_axis_tx1_tdata), // output wire [63 : 0] m_axis_tdata
  .m_axis_tkeep        (m_axis_tx1_tkeep), // output wire [7 : 0] m_axis_tkeep
  .m_axis_tlast        (m_axis_tx1_tlast), // output wire m_axis_tlast
  .m_axis_tuser        (m_axis_tx1_tuser), // output wire [0 : 0] m_axis_tuser
  .axis_data_count     (),        // output wire [31 : 0] axis_data_count
  .axis_wr_data_count  (),  // output wire [31 : 0] axis_wr_data_count
  .axis_rd_data_count  ()  // output wire [31 : 0] axis_rd_data_count
);

/*
 * DEBUG
 */


ila_0 inst_ila (
	.clk     (clk156), // input wire clk
	.probe0  ({ // 256pin
		//126'd0          ,
		in_key[95:0]    ,//96
		rx0_ip_proto     ,// 8
		rx1_ip_proto     ,// 8
		rx1_icmp_type    ,// 8
		rx1_icmp_code    ,// 8
		in_valid        ,// 1
		rx_cnt0          ,//10
		rx_cnt1          ,//10
		filter_block    ,// 1
		suspect_mode    ,// 1
		filter_mode     ,// 1
		db_op            // 4
	}) // input wire [75:0] probe0
);


endmodule

