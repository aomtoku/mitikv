`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KjBO0tzHYKmFz+A6rqum84g+M5WFU0kFm4+9K8LdlsLYzV0nngEL4jep524QSuXSoSvZyB9EUMwc
kTLH5ij1pw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
edJqp/g900AsxfZU2BonoTWahObkFSINUtQ27mA19DFwQgOzeKWKReLqpKmVUqGeZPvfHC9/kaKP
tKQcjwtRT8veKjMbit3dubyXZrylnJZlMF68gkZsNKIFGCsJmH5O//nXHmBxeIcX1VAKR8Kr9bzb
9kr0dXKII8B7kkypmzE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
prrmYtH0mJsOZvaKbY12+aE82amXdifq/PlZhaKoSzNg9RAatFfMv7wDlt/fpLNtv9Qey7tbMUl8
MkDCxdbH+Rwcuw9sPCvyLMoIiUOAIuIeJrdLqqd1RbvedqMyDzRwwAnGOASLWmnlguCWzS2Pnwvz
vGnbtuhDQTnW885p44jjGwH+MlD3UjnmN6CykUPvxFZ7FcszS4WDhWNmpeU9LlxdsauS1Vyo+gFw
dajhEELJZAapvwZezOLsB6feUnatwWO9pIMPcuNpptKclbsp0+TZ2ROuJSLXF43lqIbjOCraKj/8
mHdQf7oU45lg/R0U4r49d8BbgiC4QUMXbm+tiA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
34obdx+3WX6Rhrd9YL0JFfGkdbdojfRJDEPdW0F3Bzwx0aCtsjTdFFmk6CbLjcBqkXZ5kVy3bitG
rkvVRX1d+lPY/2+8PXXoT0o0YpuNnDJMqJt+Xf2iJXQCsFP9O72dJrOGd91dLvEPOV+THlGs70r1
CelnPAGIWlubtMMOZUo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oE480r4SQjTvFUus7cCDxBRnypFQ6MKCoEgb64GS7nGOqBgyV1LfA9vPQiVjLMOST35nGj0/ddYR
Ta4Z5X4pv+g7OyjJKH7xVhZVw+61bRvj7bDTydwIqgcbS79OoXN0TTdu80hawRESaD+O4cgSYjut
ALGVTde4Cp43wt2hLAT/bFPswr/eg0WAz/HjBD++Qmm4YsMHgONAfiju0DQlW7fpeymHCO1Ucb9l
eF7FW/G/eecgeJtWYVFj31mkp8SqVP3D9Ehn29JKNJiUCBNy1/QohdeydCjuKIKSiEyunFLfh/KE
M9k+4O21klg75W/snJBQbtyW/SAh07cdxEPcbA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GSEQ+2k94SIzE8jZjjqbUn6zyZIVVMMPEXurn3kNUQzj9WZDEimOrNj9B2Y6rDGB5BYSCwrhIRaN
TXlaMBSuD6q16zpjPsERo72vwghPswLGmq8Ffa0BgTi/w3fStsI0TGJGtmWG4CejBXcIA5dbVdPt
DwwS0V18GxyX5P+UHGftIj+lhSH99agN6FoYNq7SiFqqze6UZv4zRHmwGSduFeiz7q4qvSd/+1fk
nOYi+qUnIcESfQGzoqIycVnspHzkQK1D2JFDedglr2VHstfkd7CeLLyIAZH6oom1FXiubsrGX57h
lJeyCfY2lEYMfqt9MPl2wormDmNt42dS7z+pKA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 544336)
`protect data_block
hQ3CT7HOkkrGdFbh0TSqSPP4QaYKrssR0CAcxcoIsRQf0c4tEdltzvDmFeaS+OGodzTw6OlTWlLc
SrURhQp3an8DxBxdYaQsG22q8klukIjRZDrSP2gf2JBJ3wf5ce9eqUT3MC5V8hCZg6IvNInTu6a2
/Kr+MCuV8pROgJ0yWH4wNkvjgTZdRUeh0+WdrVvLrlHeAxU4iNid1R9BeuVhfF41INrUOH40KZKc
FgPjc2DEgLpHUrxU6ZEP+J5Rh7/GdpEubB52zyuMica/H93WqmIz2tvgS7xXLyYchAxE3xLbFbe/
SczpsJDcRuETpQgIV2VnDl8z8BhN/MriUGQM+jtNZyFFeH6DGQDraZsLcdDRPSfomGWpBnxKCcN0
SMtv/zh4EEfohGdmC8sEcDbDMHUQ8o7P/NhrSeGjrEEkWvs8FfDq8uzMnY4BmNK9Ow8pjw/bwtWy
kg+uEa1cWRvoh/3OSxv8yIiTNvRqHQ7sp3FITv+Z5LQimxzHX2R0T8EnSoj53+Pw5wlEejVvcUYh
SfL7jtQuhxXQlC2Z+U7oWrb5KZoCUgL8JIxLLMDomJPh8rkcile5lS3ZRPbzdXZbvCxNiTYbAYoM
DD97syTViLDFaWpjkvF3qZQY6oGYiBte2Eqh8km76oJAHQJ+3hnsjl+BNLIAc6G7YJkyjMY7qohk
M4QlD3ZG0jpf3rKbfsslNJ0wAPbpbmHKxyk115Cx2d8e7jj/urroFYIyVQZDz33xK8xKmz4diMRG
UaQsN2gyjGUx+i5RrEllk1FuBwtFHDQ7DGKTeiIfTETGVlZvw8nL3tZcg7M7cstf1qybeGxjcQhY
hJ+N4+HSZ8x7L71xmgl4+MYVAvaMmEXiFg18zpXQAilyN81SQcFyffjE1Z+xxe56fcBIF1Ys03FH
hnb9WsY0Q/RpTGQe9BMlZQO9vMsBoQiE4CCiR5ky2Q9dO0PakQpGghDSDvcvBtIRIHWFsaDDP0sZ
shy6sr/RvFtsoi6r++BVsrPiG6fuxerTVkTXyTuilo8aydm4W9UuHFj1q9QGlOS15ujG2miAAB03
VM41n8g3AlasJ2CwsKHVQX0L04ThYWIGKueiaCcEdeUvrB61NiP3Yguj88A5sDrrHb+21Hm4qAdu
hlB7nAo8JndFqTmkRR+13GprwAXuqo8x5bbAyz8wxK6WSiXG7zZNGhBUMowYdi0PBMRIwJ1vme6+
LWC7tSIWMrL3vcgDpYiMYDWkjtYRETFzLaiy91LfNpHKRYcc6BvyD9ptfzXIAK6RWcfk8SWomB2v
/musxjFwKKgS2PVIMz6Uu2DTFrI53/BpS6YUJxhLxDw61eCUKAreHFaI5n97bOa3w/o3kD/cTXK8
UJT5DP9mCYTPodlaUXDrpDoyH1gSFfpZIQcpNAOSEYUG/OUUlZDVrmLdq4qTf3SK6E1VA3RcZMJV
00SgBvU/1QmvTGdNJQ/O7kPuioyGg6d7AXPDWUS+BkOdRx6l2tLJRX33Rri391hDPg26DR5LOd9A
tL5H0ptsRdUwLj92owxDtHLK5fvO1W4c8dsS/GLxRirOdXBFAR9VkXh5n6eISsjWm2VgojYWPhvJ
76Mc6e2nvU1e3kErhT8hspJfvE+Jhz7rmHMO9vo12glsIqP+rA9lz45e1wM8U5hzMzSe/eluNG0S
/F+FvRM4ZIUvdvYYdTJCQ/1QFvuofu8piwz5jfVXkrvwdS2RG3qKliVmxAnUAvbkdkIKRypDxwR3
h65L4yzy0j6TWwr0i1gzGed7Y8UdT7Sa9jFpgZRTKOz0nhu/DHH032eSocZ9g+/Tf8StPC0fqAYw
xFuctVXeH7EcejEHAZeX0Jf51Yhf/vePbF/fYSz59nm2yoY0GxIbkxa/7f3ZNJun1f/0hI49bPyQ
W401Sq7VL9EZQLOv1iQoh7uh9Fa6uIFKDtULNw4MlGCEV+TVPAQonNDLqpFIwg4Xt0mk6J6UkZRR
yAA0J44IEYOUKM7LRNYJFoIonJ9uSbzVWQFxw1j1QVKCKctZSYsLsRQVpKubYnp62LGG/7+37B61
m3hOdiH52vwLX7HYAoJ4qvzGy3Yvp3lyc+sKtKp1owJr5ATaISysugZhLZIzq4XOo5tlwDeZFSi9
+2QFrcbtOKmVCfjSlciJwzS+/gU2jtmzABcXichEG4GhfY3bxp6jSAweinEK9ljl982d0/AzWLQB
Xvs4RIf/57ngTMCsRJBJNSHw4P7U+hr+ggd4jrqucGqqBq3fPXp2Nr9H39L93H7+UsngJ8HKuTAH
7roxqP0b2U91qDm5mnOKLfcutxSp73zOVCzwkyAheTdjDkBtVynXKyATjRD3WvjKn83T+/xb6FWY
utZIgRChpJrP91jkoNZCZrOwWVBI3wGd1RfBWgUG/ttxVx0zkhD1LRasKGknBT54oM000LOtd5Wh
yIp6aFCZpC+keLL4oCDEWgBvObhZiRo/PXu7etmVaiCK/d2Y+eJgAqmNbbnl7QzGOqc8Hf/HAT3b
30gb3KJ727O2LhiSyjknyUCe3Jd7GwWTQRrtyAe3fa/USnovTePKRgxGSBGRYm23enh20cCXFFHC
bHZVvIPOnDOZQb8u0qJqdg6Ev2EQslP7EyQ+/g2HL/Tp3AkPi0FiDC5T1iw+FJnfNzt9+hmAZpkL
36OZPzx+y172b78n99OaZzzIA6nubGxLoYWs9rKPAe68ElRSP3xazSxt/8y4w6kkCTanJfixPlHk
HVufnSNx8nEx1w6GRJuIKzVH34UvSNtvAIwoOBVX0hvf1USmiF2HeZsNjaZh7u3IiDjqk2xi5uHn
EUg8ExZZPMs1LGO8Jah94Mu/0pWP4yYbq0/GhjAvlg4E5ULtHnV37HUSe0aeTHPJrAYchpIIgQ6z
0BxY4a7HgI3g9NpFfr30xoTwhj9geLxmpurr68Rg0X4je/Us03yy7tp9oKYSOLs565aRERRp6zLT
9MEaX6AwdXzB0i04tfc2yVMJFTMBKDt3tRRbH3OwZdtCJRLU69Mlieh7yvn4LnWzUE7V1pmYdnc0
F/zpQ0uMs1U8kKrbDLKuag1ycQEw73mp08+Pr4mynRvgH4asDKxxhVPmPzCPJ60oWDKcD2UKzdC7
4xKnSqEb24bOB/hiYPimdHT0Mgca6DjsdxMPFNFAON5HcsCaq28xv4TM95Yi+307RGSOupp+EV/5
rYYX7JjcFS83XQJAY745WkV+8yHIdiIkDhQjX4vBHkekbx50+MeG875jTnrljA3m1Fwy2dG8ilhS
XLf8Q5jG6TGuBOEcX4ycxoRUjTuX7vo/kDuCkKZrBxiV2AvhwA29fHpHVEQRiIeDqOFpQPCIh433
TGrUFuq2MinL9CMkpGXYiuSYvPEjwoCMfOIcLegep7wZpLC4R/wF/qxQTvnuZ6CbsPNHbczCE98V
DhQ4B20mY+B3alkraA/a2LRUWi/P+DIgLcZBv5VsKnSmX1Sem9jdqk7N3JwQVFVowCqqOEBBFUsF
Hb7YRfUTlR5eM1pSDuisDUTmHyI94P8ZjLfABlWUzhJGMkPRpcYadpS2+mKt/D9OQ+u74yxA+4ic
sq5iQozm2ugcrDDTQxdbt+ydtTKlTUS+glk99KmOJRXxFTduYPDp4t1sCeC+wdX57lONdAMAhxJn
zmQYMHRaqlinsxPYgd3NrtPWFWuRnN1FS2uC1lRvF9TCLhWTp1wOlyVNx1v69RIbFA/KNwLQh6of
ozsvbauMRrR2bDmv3oAVkriqeL2tsXgYC3uJ4cVqPw49Q49vBFBSuQSGwYogDBvB80bCvnATcZTw
PrVmcgPvNKgDMsHQYkMo+VpiVTm47krhjS8oTvSr00O7e4vntLAToU5e9t5C0f5bPMTtsv7gqm9I
a7774//rjyPB8MMvPe8uw8Ew6oZVc8iWgLYEBeZikP+uCjhe+dWTp7E+NIuAkjCEPiskNQOm404r
HEqi4+L2X+wCizJB1HEKHFU1hNYDQpKLZMtdpzQKW4jmEj/DnaSQrGvGxZTA77JmH9Te5uB4EKbr
a2t3w8JtnpfIiYzVmyiip81wJhZrJsPSVxF+sDy97IO8k0intfZhETVWNoP0ZXKIwmCjYD61y2PQ
vl69Ub3eoTGG/ByVYXO2iID2yDAbmW5WLyF574ped1NBEby+Y0WrFiA/LOCGLcnr5aRWIpiSdG8p
Zh6es5HOF7H0gGUrxlWWrO1rCqWG9AJzWbGcvq0slOS/sRpB/PgSEi/okf85l9MOl88YcnguN7S1
HepzgmrbCzk5DdXolLXcJzON7SZjdlprUS74MIn8QcqOilernRWF4cICHBr0RcIYZmeQlxF1L97v
GK2EhqhnSB1k+goCbetU7ogc571A7axJm5kYPxD2qWvFA6YDRVvmhWBYxPLJ3v1uo5Kk3jyQ1suy
aGuEgnOVvehwn0cT0CBK5W6YvwVP8uAwWwYElyW4q8hyd0BYC20vf6XOKHMS+nxEF2XqKwj2eCmq
21GsvR4edGcWbkCjYCYyvvxpp3qyC1vlibldt+ywPPyMKGDyiS3R/mxgVal3MSfjFXEND28OkgdV
fHQnDGQZ8ZfQ9Pod12R7PZryfPBhumq3vqX3XZDmmrFxi4ygw8bukUETyy+JJqtZ3/MI7341yuCt
zQrE4GIcUN+8G/3VxaZsN12BgmCcjAZ7Dx+foog1G2/4y+rWBiJjPsxBeCdhHAXykrei/r+dYNsa
RBYd56krShRBVAOBYEI5ITPUFO37KH7+6M/lFsknnLP1G+MUup/i4/arYaXUP0jNl1HlGL2LUinb
IFAs7GaIJ1aSl+5HgXSWO13SJmhXkhXxH5G4gwxgsr59Ep38q9ALBjgqY5CY8LK9589PaQgdatcV
F8IHGZfa9JCOIj8eYIUyhwFKxy1LxlMsLj7tnO8Kos9aN2ebHs2uRd3L68pIz8LwRIyKvmsNjlJr
de/FrR6grTtO2e9oG/ymz92pRTVA2T6PcW8h3dE9s3zBFhXnV5BgbE4NPZUIl/dNU3RCBsW4QmGL
Lyj+iI9s3K0xUi6iWAW/LjllOlKEu314/Hl/2tju5yzGFWnFPEJM5ZlYu7sWnJkng8CffkMPuVLC
bXbfpNa6/Vh9QYlVVynm6Uy4oh5aszvo64PsC4nsMDDWZpq6HdYPfT9u1FoFVouRZPYuwhtPHbW9
2tjJ+KNiqBHzMYqCYl+62uqklcFbNuj59t2XPG+eZ6Dz8OEechYQcNe8y+wgDdmt5mcpoYfwQfjI
INL9a4H97tYhNrmym1QXiVDcyGzAt3HHndH4Smjj4ftFdSlELsFDoYSEgcVwQgHFNnrVuvRLJbs1
9FrTFExdAxKfVqHw/IOmd5CM9TKzCv+Pk/lnD1+vXuWwUsksU1Za+/lJINAH3GgYktRNvzRIaRt9
RwznaKolLpA73WUfnhe1G8YKP4NTVq4V49jbQ2dRSgTYRNHDzs0Af3VvfyTy4mWcvPXYt2e+Rn9R
/FMiYph0JDNYXIDSkn8fPVkdyAdcCyKxmKjCK0EvKu5kLYBuXIdIOlySBXGa4Uze4+eHs6x+aoPX
cQxoyV+87SL/4wZggd56Uj/DiaATOcBqph2seIc3kzmSHl1GeP7nhLIjMY90IeKSlVznpuBO68AK
4aZqovvRmdaysNMfhop/LioWvMn4xe4aucxHy6BcKsTxSgU3/1MrPq2rDYO0+kL5gYd6CTj3Vt/1
/udzJpfi2bda8exxk38bBbh8EIbKmnHkbuj5NtdUHjwGiyYEHdsh8vziZZKAzfFZacLfK+sc2Xgj
9WcptePEMvH7OaoEUa9wlwNv5g6Z4i/sNIV5434zBVJoUo16dgq7yTje69+WjmcWakvwRHHd1m8b
yYvdO8VSKTi8ApXdawb8cIQ0psGQquTY7Fep1Mv/aW+vZp9mHwoGKtSIG+Kzavm5yPblgYaHbaXS
0IZpVtd+2Q9w2oswLI4ZeJNZmzcTcFPtofKPU++YR3s933GXj7/NSTssS47QTKSL9e3RwOLOp+TN
2oW+/HpYsOB4dfJ/zwTOzQxQsAoLUWIcrg5DAkoNk43zvLn8KpGrG6A7E/MJ/l1VFI2XlvJrb4bT
vRDs4fd8gYFLH1sPfs/ITvPbrFnjz/nGpHS95VwMHI+MMQs74aJJ+X4zUrDcSEz1EHuoIcde8Pbf
qjPMOf0yS0vTD1Oy80BV3VITf4dYKI7HsOODndc8tbew97CaSiWZAnOACATC7VwWKFkk4diGanCB
IyqbnUM/FrNU0aw3pqap2QCxfZqZwmangnbf/ro4OLAULWkmkCZXReE+E668YyiO2R6UFL/Vlh9H
dMvRvTXzk3GTUEBG2FDaSlVG/UH4kR/PGwXKG3YP9t2NzVkw1fwiAwtsk8frEJqvbny/1L928r+p
eAOnyxNS+gcftrUfB5b3QpKXtljnXOlrQL+++UDd7orF7T6beQ65oMLpH3kmg7DxPttMvWtt+OrH
XfFRvENCdiCV3dn9GvB8zPI+j/Vyw6rsKQjSQJUpsZ7p9irmSWMYdgK+QJJKgsELfWI6iVOtZss1
hOZNK7tqQv8k3+SyS3awqfpTvGTVrBX4MuIazTOKXQWZb9FRfw8GnJLczG76yYMgRiwoaFLMj5vi
CLRqGNkFvQyjcqnhlmdn1MPhEMHf6KwC8f+bj3UFMCscycqdYoeWZ1OmKnm4qC9//o8igoYQ+Eth
4+88prBF/ZtK+0PAaeI+3I+UJlj+5WfrBn/q5oUTBaHF6g4/xD1GHTmjKRpUkusHsH2Qtr25jB3C
noa/SojGGqLc+3e6wmTKTLw0DNvCyq4RO42p3cOrvW82kOEHEipm+q0y2bbWvmOZYjPP/Vlra6wD
R4p+iTlEwCUcGrjQ+kzKK8B3TtCz1ndksMzkUYFvIX8hsDi1SCmR0YxqrE+JeoZM+iFjCyFWBA87
1pLtQGD0CLeSVN3DxqVVGKGh3sn1USI7vaxAlCkLDV0bP+9n1y2IAgqtUeb5eTHVUvK/gieB5dNB
uwEwbaifW4eW4OJXwOA0+zaK3Fw2yNunegRVSnwSQSDgOk675q182VyQxt75nRNoNrk5RBxxsLel
7KMrlT1HV86h42mgS3X4xGE0HEAURKv8UiNVXE8EYCkGJcUSPHLqQgU+z+TOUQAg23oYKPPKYeZ0
nvR/EAdMNn6E5kRZa4J/2pbFDOYvnW7l4/gKJfvULaHeoTjhLr5HXeBT3LpUiJxG/77pSQ0vSZ7v
wthw0zkilpyPiiKrE61R0/uR2/ErP2SQg5q+XhGfkMdSNQ8HXSH5trXSVD0anwMbG+sR6YUhGSfn
wyahMfWonBPNPBZ3zvhvOpdh90BLIAIgO+59xli93v22rQKrHgm/2u+70AqBw7Xoz2PUlVMlAlOA
SGwW2ntC7kGqi4BGkyKnn1WalVAGPmGmh3GY3hXo2dzZ9YuqyX4bG6MY/s7ZkAIF+LRXL8E7j5rY
e4s+LhHblEdJabGhNkdY3s4X73cQLAF1PBsyVDI8yDzpP18PYs10+jCnMLUcKFTe65xDEhJWi8AA
LZhvy5TbGmJwsg+83Sb0e10albVPL7zzOuUhfNP/0aC/4k3+jYR5g1ENjGYP7Oe1w5kdgCKG+82F
rjxVpZYCoYW64dp7F1eNCrhLsb6wx93D7PPIr6+vbmbe+eDPourAJffXTVbkVCLu/xc8++3G9eG0
5p7Jt8yRz2MUX1Q5GUmlLFP0Px4oN4iheT+pVb4Y6HqTBjArpNjwtk1ruZ5sG0TOGPwC4Jquac/u
3kglEfaR4dpvb3AiUkmBmETIo004wpjIFQnFdAwjQ07Px+7tzyfSEIBE1Ma6N6v0UvdVDxZTs+bX
OZaq17uT8z+tVgPwjOVJbzWwJI9HRZRkpZekSrYohRPLH9L1S6Jay9B+VCLoay3CyKiqQARZAY6a
tH0T6FOQww7ky+zV9j0w7MOD1mSIOg1z0Fo2tLScLPNzNCWJO5xRGHP8YdxdBYO7fR/Z7YzrByao
7TumBtFPvgr3otKQU2gUP+8Wyk2YGlTTFd+CkOJTZrrq1693OtzRD0hDDjhuGHIW6/SVdFinMwOH
0sS37sSRVOMwraST+SyXXwuHHOCrCa/gxyZoI7aP2pcidyucBioEN3A4ipuzmpRsU1leTn58ceIY
IAHjv4J5HA/77Tt5oIFL3JqsB8zQLk/AcpLELG9/2Naim36UCnK3UUCWApHp5FIcDpsOyNudFHMD
mt446WQ7Np/G/aSgwZtQzFjBJiLsLJCfBeTck2ThDNH3AL3QReJgVXjEYIUm9f6HTFqCC0wSHUjP
Se4Kv7SkM7pMRXZug5+L41qk/z50wD7BPE0qD8ITwvnGG1EL5EbVp2jJ78OxF1OlmbVQgNiRoThs
M//YbyWJUODQdJP317zhWRkm43BpwfO2tvQRzrzseLn5sNu+r6bfa5qOQtQgvNjyEhM3SjaR2n0k
mRjXOVWymnaiWmMKPiFG8sac0T3XZBLI+dUkN+lgSrHl6TTYq2Mk1PeDoRJbeityKlbfyBcrCuyQ
rfkbfXHOuyc8YsbTgRTO+/T8i5dAQxX/fUVqj7zsjzQhMaMfVxS6Rt72D0PeU1xlWQSKYLr9mDCL
cI24xaWNB6RhWs+KbuMZbGMViIKeOlD4JwqlxjliytGU0UyfDuXrGstwZrdTMkSQhCNWgZ/D+rMs
y0hNEfcB0CzLplMAPr3S9I3+TqDzt3tpNX4yBfBsR0pbBSlWku4JweKBvgRqxeK2L70pecR0eCdz
7+GATL7IDi9hoogbbjrLY8jTS2Hfz9MymGA0gjn1/lrk+VwAvKXcud4gfUy6QN/r6qqapzkjynH0
p4jXPtlL/u3WVbVcob9t7GTDR+EMsQEn5seOpwQgID8U4fpZ1omt59HZcHDNtQKQ4sYzzelXpLVT
9sm6GRM1eDZuPq8KMKDjOnFQ2VTjH7wP5CnN73HX80zRCuCnZj9mgHOS0KoHy4NUabUpVwgF0MUb
tpy3UrxQcsmO4imeHE2PuH1qdkD7RL+nqXr9c+2Rcp70E+oYi2sVpJPgzNTBfBG+4ikPO2xE0Ld2
29LF7S0LE5hZ5I46ZJmUt3lN2RgHrobRcsgK5dIxKpBeDd/Osa59A7dB31JMS1i8GuxO19H6FHwc
dzhUxGNY1CXzbRMsiGeX8VYtsE3/9+mloqt2sYW40VqmuUxy+N9FEftlYk6t4VnTupzKGd4v4JRP
+9prJo8JQp1iMrMxvpq+rEncN8iHdGwIbwM4Wm7IiWFjZGNFhftg0W5RaWxoYy4gLpKNDPkMLow7
nXRRMZqiBS8WKTbwi51WBGKFnWOzkhsVTHxmsl1GakDKqUGTYusOcRELa4rhHP4td4Km4iJESR4c
rPZpXKTut4xBlZQ9/Yti8WpsmpB00uEq9dFOIrgUXtdfors3arVONZuozzDghkVJt08KyM9SYQpC
1ls2uWo6QhptofFu5gS5h5Lw0R4YanYBMwdFswENrCRSP6447xA2kT/1VDIa/S3MMm+uv4Hl0SDg
Wbt5jY55eFnieuRxASWXRkyEf7ZN8L6m5q+HzQhJM/MyrFHeQxonbgAq8NBBT8Y0bJDYxKR2vUmn
/CugIh4Tj5Nri5/YYguBRCecb+2JYgnT/WeTnG9DMveNm0kck/+1giA/SfTpoXQKknfGG0q4SQmC
7VimVLZ6H60S/XtcaKUFg/vANbcPDbhCxfaknKHH+xR3MuamfPBxxXHovp31r+kAw+qT+7X70xAF
Zw3426zXr2cc+FADNMP+zsng35QXwI/uaKg/2wpHdDTL8o70BRAnMdmSW5KpNnj7n3gFY1ibKejR
MqRcbaXRpnp+m5uyfZ+On/x6tf1g7X8A1RI8M3Nvja5It+w8tvtqLTjojOrqviKGugz+lYXFBZIk
tRPIerMPutjHNYv8MwiWAzO8vHzwj3dVHqCQnmzMsM2Or0GZGaFSIg09aODWvX/mUVDfLVINvhdC
vi+QLIjMYbt2ajP5yu3fwgoi/ljZ2L83PkEMZPsYB7V5HeXu0+nEBwXz26YSTC0h5nve8+W7EpAr
Aj8tausdCufiOjjx2yIigfSc6yq9ihr42xrxwJbZXx/icXcNwgJFuMRqRrZcV43vVSdK4ix03wbv
qH1Js+JmNyL/RzhHs9uba4a3iMT3tp5bCI6Bw8jV4TbuTij5yBhadZg27phrArnBulmM1rYLXh/1
FueEBM9g5fmx2xkJrNKCo8skPNjApFMYs53vuS2ReUgT3U6sY4QJ9c3f8bwKfTIyIQ8d/MMMwBU8
f4CFNNfeHcLx95+SXpm+gHSh5D2chCnTcVtTL7qCcpyWQ6LMp/TL2H5Pv+yZfk7nbKBJK5L+I5LU
zW0UKfekucaAAm8ydIyta3Vrqezyx3Vz5FCVR06q4Z85+5FX0rMvUdERV7ecrO5+M4HjFikzm1HG
MtcVsAR6XmviZIvEf7Hsg06krpnbCGsEpvflS5w6xxvi8sx/ejHL4DjoYR4zLx6Of6N9cSGBwNKM
K54EPLDR/d5lWMLLcLW6YxImac5eTPOW1hY6s5BqCOeC4Wq7oDLDIzS69b7Z35s+d2NKeGq2jPh1
/i/SONDQHCo/eF8pM92DHPn4DAaAyXSvisYrvdLB1uFlSzY2F1eqN0ASXGCGCymPZ/5gurVzvcWi
df7WO04amfH4cxf3X54HHW+mGnXxHlkqQ61EP9c7ekYY5NKvf68t0Ft2yN44kaAEDqKO5+b7i5wv
lrpKlz4HSkARI9/JKpmsQK8Zfyg6T5L0XP1863D7Gnd9Fzx7Irdd//TNDaGnDGJjl7JySl0x7xFm
+eeXxOjokonb0+NfsqEEUd7ir/Inezk4pa3aAvEaQXqXwN5LapAUEIFLpLohA+Aqh/WyIbcTH3Ts
LAKStVSMFS7w6eoMtQZ8CsgfsnM8xzXMQWrEuaDN4sJaQbtIKi0m37pYOo3B/sWPHBhOFGkmM74E
Z4ENpee3ZBOzc2Uft0/sSkLAO4Xqfjf3/jAjnL8FVeZ+Jg4oEzWSHc7fYfc2RcwfV2krcHLn/P5a
6tuVBK7VBV+g7CDx0leqFpslSBYpO5OwPbQqHZzxd3S6vNn7ukrqBq67VmxRF+GjjdJe53S66qoN
08MB81his4OyIxuVVi5zNlVqQannPOREkQ4P/XfyZCW5PDtvC9OwmJUGIoFYcRfT83Uqngntojw1
HQnq/qnKfaSwS3p60bPksE3DBjZzGo5UkzgqcqY5SjZqN/8kDnizSbPrDoJYDXiVDp+5a0xuwyLD
99ItVq2YUafuZ2jV1jnQh78luQhs+BKlSQ/auTwOS583LcdWxmxRIsakKIze5AE9ruliRozN/hFX
uvkE2UzOI3DCWyUPK8/ODrSBwQ+Cd+tFwfwcROZ+yZbXzRhj6dB0Q7u30Vq+25Os6SwCbT83aOZl
jlel30KoPXHU9to+w+v7YWqnHH8AEsTf22itpIWX2SJxSszvApETLlmjXvOZEKeSn7WHXve832CS
XKquGgc2vceQgo7fJ3HIXYmkfgqiCXoA9YyGNKc9TvvQtAlXpAf9JzrJh/RcNv1Fyc46g+nytAgK
Lfp5pshsX+lmRT4c5V8sJJL2Ebu3wrMA5+z6NVQwo6BUTm3QO2ycy4u7GzODWxd8HLU/F1NaJO6s
vUg5D2R4MhfPajNy3wekOmnuoDSeoahiqQdklAXChxXbuSjgnGW+PI8T/hW3VgOd4DBFBJ72f9R3
zQdz3ar6unvAUhGrl5Vdyhck3/9ASmCtmLHMwFRNVnmIqcPiX/ooSZMch8iqNtwW+NMcw20hxpba
3sBkaGPqYj6jFPPMIE+UcMemAxYXdOtr5BR3UveOUpqQrO7wJ7Zxr1DZNUgfE5+f+nSNq9RwJb77
srNXzf5o3g5SJ8hrMojzrPJScnmngJJ3toe9wR5U1axhAKOU85DNoqacymdIkq/G7DEZGHQgJM55
D+CmJfVpVsAW+7sNreQMQZFaP6WFmbFTa94pYhcPD1y/owbWAJdbgGshmQU/eq31fqizJNwfo9c+
bUtS+0JqoN6QDGFkE9SB4+L9Vt7gSiTPUXY/LeSOwaAn6MK4rByPQcmSJEuoIN1InjsaUpbVWGEm
/HCFLopb0S73ocAO0eys8kEcsF67W/chDoXU+fsxMwQcHawiFMZBw7WVkwhviNn0z7T1YIpozk+g
7xgHvLkAZuP+y4GSjPCyB1jOSPrngo3E2upXjnFxi5/Jz4q2ozx2ZkSviDsNcm8ss71qhrGuqlrq
xkpYqgdA/JuxEEgL/VVmKNOhIJVmAl0cnIR2mZAptBDYPWXbReNw68spQlzYA7/ArAotO/GAdgyU
se3zpao8J/f/a8QPe0N9lIp9Iftza9mywBiv9WW24K0UjI5WqQZ/fRRk8dkgf+raV4d0JvbeUk4F
ruoHJiof00DuSDq7QGgyitJD4G/OuJnU1t2F5FMQKRN1OYCjU/78syJRhAiqb4+ac8CcNI60RGFk
7dSVUpmU7Mn7X/8HUJsqkb3+TsLBPcAlfZIegGMvsqN+eeIWDQf5bn3ulAq4jUq1/cMmN2A/xSrW
ysi3tO9kJ0KfewKG1pOK0HpcY2mTipF2iSAiVyyyGGMYGQW/aCpV1aQCO840dzLki5IhA9Mf4c/q
5YvSDfG4b51n7NbDjXlzNCRWVeML2Z6nk8Uxdl+ZbiEEKfEjQyViCOatX+GyX+UjVD3LA4rLuPEG
9kQ5j5TK6fLmgRob6hujubLuclW7vPilFdYhX1Dwtr2d0DN5cJ/MvTeSIThLRQiOxfaMxS84H6vm
bU699TWpcy3N6oyry9b64IYmir7I6retZQsWWIX3J4RVzZD3TAC73VxHE6XGxHzB2TBZ2b27Dy/6
erm6kLBDyN4tF3aaJwBbF1UGQDd74kvlO7TrZIy/3sfs4pHgHiTSuEfaHGTM/SMeDW6gTWotU7Ky
nQy7P4KyDojwhRmypTCfNSGuqirKDg6J/2nsQ2ip3OCUkLIhF+/FAQA0sO+Nwsfb0uJk/yVGiKCC
HcKl6ipD2dxyWqBhrbeWoGvjW5e8BYcX7XLInbAQIRRfeZHMSUx6PK3kQ04PBRVpS4a6LJw9X+rJ
L3VjOi/y9uKwO2Vsw+szzzsBjy+ZrFlvZYuSYp8hagVQUPotFbQHw8HEjhxHyvNFnkicrgWnOK9r
nXvcjoaZc5LSr2dss1UMtcFGjNVOWxA0GZVnG+gLa+yHBLBQFvdrsn+5kKIJyHD6MWp+0/aXMmV7
WUezAdqC12qOr7MBwnrkfCjTFi3DQN+QZMF+LyDrJHt2Sjo/sWcwAa7rcp2T12L+vunJ6PAv5kDH
/UrPngfaFwW5at925gzONcSoRAwmc0owCPRUe4nlwiqqtT3pUsixdNX+zjhvsor8jpOPkXWWgD5V
4sni/qk3mzBLm5dJvahLpbaGUWx6SPwRwRn9tvWFjA55m/INjYWYa+FeHCd3l6bxbG7qHqQHcqyF
f8tngCO7NNaLtmshOma/eM3Rj1KW3X8NFsVP4PJ0vrkWa/hfqpOJ5evqV17NxaU/6sp1GhQnmr3e
fKS3yR8l/X/3xO1BHM8HTE7+nMu10VtFS0Oaqliv0DGLYYXIKXunp8c923KufTLO4hqdEJHCL7aR
Qb1lFdJw4vsP5lb1MVV0hAoRvPeoAehf+5BOGfNEaJaXsZGLf3sUmmssAtLIoe+DtUuZ1RcLvsAN
p6ZNuPCGBSmCArWFZHGXutnZUIZLUsxt5DdcHxPXxbWFGkC12biApOU6oG9ae+uNBo9CinzQOlbB
EjZuiOkUUcWFaaO2igIwhURb3KdhOIqCmEp2B7AwFn9dEvT/2t539CD6bM0PrIzxDjPwEPsSAt6q
x4G42kEickXFgOpA3x/BhrJ52szYgvmCH4x2SafGeB3T1YyxXU0TkTPpqEAXRkuz3ufIkwxJM+z5
nbpvMBG0l0G8tQ4LgyxSjWYr/XK3Hp7kLwkrUPOrZImRkFQNtwniFck8O/iRgz+Yq/IZxOFeyzpI
qZYX7/JrTYJv6164X09/eHp2Gy3xsBkfJPbpBiVWQEowuDfsWU8B/Jywe43c9qEVeEynvRGJb8E2
zb18tQjNVgKjynEcYJIOutb1AHqMd1XIc3QcR85jwTdmxMNXqiydpcaGBxNdCybdYGExRDqwbWgz
eym93TGC7u/5UYvi97/t/W2ZFhFeeTbpoEGTRXHO/NHx6yfi8IVlZoXp/ve5rSUmWL99tk9+DAxE
YvLjTpJp+FtZzflTt3Y8aWnXuNruY8CmBO+4tvgEm9rfIpbTCAVnoGLbLK7RC7b9iMH/GSBc/8Jy
hYzmwfv/NRbsGPXKycCZqOiMJ2vs22YZHytEEoIYC959SUorEPvAcW4DL3C60OcPqEchyxmezse1
i6eyQl77IEYr7EkhEXdZa887dV7xTVW5LWX7As080hSmoHGZLoTUgOwT1reen9iT9BO4+FV1c3sf
XcLWt1iaNtLz2Gb0aCeOHSM/jJkE9I73C98UuWmAhR8ilOauquR6pVawRAjzkeFxlOnJ0AXDTpr7
oJPD+D4TaPibZWH666faenNt8ZtOgBluf3HOVWJKtbIzqqhrqAQfYZ8b+SG3k66u2OFRj+nr/8HI
ywrRBPOujVx1j/AjZ14BGjDF8RQzbv4ctyhZyi4ZnpY2jC/TmpwaT4q7UhHLrrmukf7i8vwsYr1U
DRiJFdeNfU2IZz9UV5duEZmUP7TyuRDxk97HxKHU+ZPFiFANr2Vy+7/cPuumdwMeyy/IlfrJyuQo
DHybilPLyvCL2DFmKs0VQZFq125DlCfNDQmxFEklwfxj9yJwqjL1QNAbdqVIbKMp3yXJU4R6AXvL
smmxLynTT6qj+c749vP7tbJSWlq+KcIryYo4A/th1k1GpDjQHrvBCwYa3I9IsscXT8hAMtA/DWyy
O13zAOQtc7xFha/CenlO6KR04LHFDmPQFZR2QUrqj+2y+hBi89GjlTLhJhoHfy7Snv5lEcwIqVaS
K9IZ6EfSuJdCJg2e6WFNgUR3R7MV49ogqWX6/9F2oGdsZOlZFpbQhRncw0yUbUncb2LJeBzK47SX
fy8BiHKOOlw6XjB3j6jmMMmwM9Bz3Gl93WODSq7NO4qC/aycaSyqjBF05k3pvcEoHrbQVAQp22Eo
BDaYvh5F4DLl9nk5m6kizfVPExH2/pKcpSBvJ+QnYY0i/O/aHWCG+1p7Xz6vvKX4r1ZP+Q/r+H4x
foI4gcUPW4ZjkIxk450yAd/8jTBG8J4uFtEdvPSkcvZzDYfYPByIZ0vi+xblDIcEG+k7orZUfMMJ
mYXpV6KhVrex/vtMK2llWf0jINtx6FpaZ0hrOKmtUGGRNxWYtZ3U2WtQXqRh525cqeNIIny7Yxqh
vpuom043zQZPrkGa4u/2qvZPqZdI6oOBKz1CbUm2Jf2XXjbGeP94RxEcJBzy971qjlNhFKt85FPE
zTIGqIMDHE4NU9z06ejG8nDoCcDWT2VWSMXhAYHw+ly8MzHRZz5eiUT9+VpaBDt6PKvUbWceTR9l
4al+pB62RnnkxKyoF+hzjZWFd7qb+wKiH4Wg1tjtWAZg7Y5dJ3c+fbx8xYTBdNH9RB/Q7djHS3m5
8fVBJtyRA7wAomdgPlfePRDr9hNZ5J0UNtUFUS4QOZeIqK4m0utIagHSdGV7nByA/xIVcKUemEMe
oUtaVzM9wO6uLIp01UNjwvmnU+RjxVPy0IQJC2HdE8C8Nu5hzNfHAmDi+ZSFMRACwKAy6XmF0xXA
hnwI9uxvRCGHSQroN7NKlxjJAKmUhCTInHa4td4cEqm2XqBZP32nvVOUr5vO+iZnZ35vFU0lmszE
SmHqoVCiRYHPEGNHQDVZf/QJNIwUBUfAWRu5aqgRTMmxZhOWznI1d1FvsVAqOa29nnYy2EUshw22
+n4VjCiknm1ZM5gVZfd4kdmp+msj7ZflbdsqzGhMqP5LMwLUndC2FiqAzApZgnIww49U9hZlwRQP
8AOgt/CnCNc7KuWe7SyTK4HLhyrLnEA+DV1tQtIhw2W7nGn3ecsiAUZ8Yb98W7WwqTAZVMXxZQX9
qi4WpmLgGHXtm6yWeaqiIT01Sdh+1c+QPOVoW0Q/Yk34svwp1EIfBbXSw6rhZ6gfGcSIw51gEhHo
4wyRpNbzGrD7oQkGXd77ak6hMRR906RPXUxbGfih2+e5xs6ZwHl3O4rrgwMR+OoYwnhq8RjFvXWW
B/AZ7oYt+gU6jTGsezQF6HbIlKyaVX25lrNOiOB0xk0yuBpaA8pfxmDSf6SezB+gt1q5HVPOKFvB
gDr5IY7QGM4/xoEKns1g0WCE1akmoC3engyrZ+RxBdDqztfu0uJI17HpjefYtsmTPP/+dTUH5WMB
/fhavHci+rODWjz/8pOd6lZ25m9DbntbksLZSeTO0r5GsdyBRfl17M+X2hqflOaDQjiHQGzepTts
5+Ruwgq+tuIG0VFj3sm2k/+F0jFCheOFAYJdjSAuCWKgHcGA239ySkX8YIWfbeivzkMn4yRCxsXx
IphljX0roOYbXT2c7roq4z8nN4XyZey56DAasKR4fFI8C99/z5h+kFvMKCeKNMm36C0jP3wS9xgI
iqCGkZfo5fKJXP8cMrI7Yd13VgcGqvocipacKku3l1MS5bjBKW/dPD5rfbE8msCL+duERe3pwAZR
Wx1JLLIweEVc6GYxOowANALLjTTzzG5Wmerly1fxDpt4LR8+vHhCBCiloAE9SoK354rFkDBBmzmg
jjWNGc1+duoNpVwIFtl9dyPZ7ZN9EG49PpKWkd5+ARA9TttEj1o8e2WXk4IWLs4nfBPSeAZFPv0p
PCVIcStnlJFWhKj0SEAHKtGZkjenVIoyNlbcwcixs3/JTBUNWCqEYjRsPZWuW+lHvvPcz4iXtTRt
k+328A4Skm1mRDsJ5Stbpq9YpM6aEo49lc5ZmhMDBETzPsFNgkj1gSweOfyu0wbvR3eVdWAyzn4x
8hgf3O5+g6pSuoDKHcEZA56yvkWczpmGFSMRP4D0SNGg03cnKDCmZgoHs8RnHn+T3zoKuvxrEKE9
Oa3Ad37guUiZBBNfumo9sPMQ8CPDhPO88eDK6wOFSmHb7lL6CJ09i3dh9HUlx9deHG4wORJd3thO
OvaARjEZhAzUSvDlBnAjabXW+kA5/vhGI//I18/zsAVVtF+kKaP/ygboWpDyyDEBZH6iRoCwig0c
l6vxV4s8tTAuIx7JkFwjhe5mr4ZI1CBfgqQR+xaMr5IhpIw2wn13S+dEKTTtAt7V10mb1rSYQPmX
aZOCNm7mJo62JPkNym7CRHXV8ESMGNxSiESgpR7mD9gxkXTjQO+e4wDwFqXcFqp8fV9+swooAfwi
gZsjdtZtlhE2GT7TOx73YjZL1H7DcQ7Em4g8vMLtQKDNBn9Y0dN1bkNHd/68C85tzPwfKL9KYd39
z1ZtFo5BvxuUcBk9QmiW2+GIf4OJcwfEhitU4fdw4F0kqe7mq0BOM3fy7JyT6YTISxnXbG5f/m0s
f4y6wDifJ6lHzckgmGmlf9KDzQPW2sVwxs1/8VyqT77hD4q4OYo7WHPDfMcX1Cntskro16cdErxH
kru7DDTFWfwf2q/CeLNpqW2kDMErmxL9UCZCYSWNNn8Vv/KWpdFxzVtv81i7eyIIiKgo3PM0PWQI
SC0O+uWq1cLp0fu2F79cfoiFNlfmPDj3WIcA9/yCNsZOUtsXs7nSzx1yFZzsySD/dwgN/PhK4OQB
/MMkXxKytEMnryIO6vcE8o9qDblz3X9DvkpCmmtkuErDHjMLDYmWhlVVbZLqEoheP6z9qGi46ADx
8701B7LRzEtKNbmUrNw3wp0N1ue8ycW5mviLKLwrdzA9F8Eb9DcIbDFJsG9YQBYkMW24DCih3A9Y
7RbqLcEA/2p5HaUy28EkeN3h9Q97tYBHPRWlv8uw4w17HOSwk1NzTucAvXE4MgkAx/fJA+wzDo68
RR1WCJ8lTU+mqt8tXGFVfgCqtu85Cd6NLV8Ehp0ZdTdKijJd02OBwjRV5F+Wh6BYm8nQxuDCEscl
RqkpFATDZyv0gkd2OZ4C/S6fCz+D4NFKde9XBz+1Gedpp0N+2c8APfOLnc2p8JnzGTtY8rXUJD46
XdOphyeY03AC2TMP+qIHnU3F1HITODhz4oFdNIgBxN5qK4wDQWS2AiuqpO33J79qvhVkb7Vg2OEl
Rx2zS+WiQOCcrkqo4DZxygtXGdBL+Tt9f6kKG3MhwHs5kaAdt/gOKGT5UMxaLvQpLk6hsSj6w6wv
kQWT6mp9Ize0oYRaXxXuqzea36yyTcfAgbLSc1p4l77XTPrh83E2saICc1OIvjb+9aHLgvqH2baE
5C7AkIddFQN6HkgDXp8QLpyH8qLoA9G1K86NIcSKnTbK0+i2WNTcpyAPKF1Kh1kn0u7QiAG2GaYx
IYi78FQBX9EvuSrdATi4tVlE0fWVrrZt7itr/KpTtli7ffA1wzdEaHiLCKsx+e5ERjNz6w5szJEC
aWCAlSJ6ZFRAiBNp65bEX+MwtI66ZaNCPJiIr8ojLw+PBn8fip6SW2dkiiIMxU2qFFGIlVBZC/QV
pQUGZ/RK5hT5Jx29QaNVuqZOfwN3HbCfd2grAHKmUvWYLwCrnmFlk5iA0ps201S5JycBQ2A6JfpW
A4mtxMB1Tk8yUEkj+6r2exXoqMOtOgPaTi+8WMT7eXhiA9KErf0YJupb6Fo9xiyE9z5skwlkTho8
ocGB18MpujyO2YxzhzQcsWzg6ATD1/5CMOYyut1OpWA/o8QjGY32uWKQJtZVCOT3PCZs7AhVLWqD
W0Q3mhHMbsGavbXv9LbnGugE2QYuxrIyU05G5SPZc9f/xO0rfoXHCBoPl/YiCHW62ojHKnVhtpGp
5IMmlPYF0uXSDoxP1g+kUL85SA1TGSlnMZOQ0l9CTfYmhFiaqmgTwsqS8ym0nftUXJH9FXmAAJIb
jsxztkGDxcUZTtWCWoErpz8x09jqsKpIXaeENYVrd/ovvJP6iGf5Z3F818dRfBAuMoIMrWHnQCIB
zfTRgMfpLOLiBuIzLRXbhCvHqcIu9MW9hpRuKZvD7GtzcI4+h6/c+KVn5cwBM9VK7yhEiK6fWH/i
RJ6N+RMw3iUiR0OGiTGoLkCRlmKEGhSdkVugNiI4UMLasHR0qtVtx44wjAoXOlXKEpydG8CGiriG
ehsz+WB0D8exEI6JpQorM4zd1bYEs7+q4r8yfanSilCDRo1YyLecLNhnEzRHlI1f44doN/nmkaZz
5nfJd8r2ZJTnUdwafoTzIjEPzEZaGkfntBY9KTCftFSMqy/zilplXc4bXRhzTIGpjNznMwwuMggv
JS8uHyrKU/Yjea3gCy1Rf2cJkH1z5Hyulz7COqgxA4/KiYp5dZ+0IS1bhLGfnePFt41VxHibypJu
onfp52ti331xWPK91mNfylChmmjkG6UaKRZRf891mzmty3RF5opHQ3hIFLGox0Oxc/tUx56eV+xt
ti5le3dbPwIKAJW3+ONSIhQOMMPvZ5FHM+bxpkmoSbpW33zyPbEVwFnT/mTRF9FaW+Jr9syzOQkh
j+ux0aNlEnroQ6xW4iLUMgdKNK2dieKGcuk82ug2XehToSQIPL3+g9r9M52jp2b2UxapSOsnF46H
xp5rj9yN8tpnUo3KYFEny47X8L4atVqZT/umGnCQYsN9snHOStmnuhDaJeIUFp34DLa3kwvEExm2
GUAMSu/zaogQcQ6xvUYPG8EeNtleEowGJuj79Zfcsr8a0+8XWN7gajU/uhVyHF5dhnjmFU7F+XHG
d97cnZQSj04jwODu3a87/vVd1gx/6swc+k13LI+KtqptdVE+yoLqnoBHRXzSpHhoe/a6dhq6xikl
OwlGgy9oJtqmKFVHiIJmx4B6Mpz8udnK9dxhmr047qwiE43Qb0agn0Hh3D9o0v/LE7aEe7pqUoKN
VmdGhbjYXb0ZOe5agBVCWrLnwUzciFlwWIZlM9PM7bCH0GjAWOqsOVeAzfGPM7WUXjHEgSpsxwxq
EbuHIoFZix0eOIE49dGv0q3fIgFzQ9xa22gnxXlSOcPRx5dHqoK7kFkvh3NaKE6fzJqz69/auTm2
NhBliQ+M/ZAmmU26DS1MH8OgX1hdWo6e0Wa72xQLh0vsIP7mnz1+1dr/PU03tPNVsFm91Xth2jP+
xDoaRclNWZz1BsjPVhf7DkXvqchqs/Y+X0UQxlp4h/deW4N3C7UcHSdCF1mMOgcJqCZwN0w5RT8T
zHfsflg/OjkwOduylfME3lo7E0LqucXaHbBq02HgUdEnfO/c2yw2JKVyzSbpvi536OUqGzSaVsJ0
HJEpWyM8NJdKsWG30DIl5G/kZL/Av0elxsL2/EFdJqWX4yla1KImnUNC82MsM0XK7vQzYgZcVKB6
EWlXK5WLWgo+eICOKcW5zaW6wQ/xTQVRNYzduVR2godtpA3MQ7hOulFQ9czIhtELYHZQDv9f96zg
sAPG9ZLhooF9Y8dsLZD/k82N33rSFDIIdeu0rFtlUlVkvcDwpr/9QISof3BuzyaIU53U6LzOy5QI
lTj+UIsx7MyG4dSFvrW3WT4v+uiep7QJMnz/A9T6pR0mVn3NvKXNQ23fdkk2lmuHsAZVcmJ7HIyu
D5/vkSKVbOUFNyZaYyO2Xv6JXNKc5FV1aCFJmnu5TERiEDGHCIjX2rgXCJ4y1mgFuHmST1l5BUvT
5Y3KTxvSyoZW2aEc6vmf9wa0Hu4/IL/VyWNqVGXmCPKjUw3yHmjdctWM804l90VPvlmmXTSKWewQ
KwdvsisIF4NEugPCYZytGsqPIjvdrb6ScDBAWWCKrdQVn60bJFLfivApb7N4GLlNB0y8xcZxmq5q
gfcj4iaHO1z/wyW7PWjNC4p9DDiN52D6xrT5KsnBTLU5xiYGhKMKVtDRHnYwaMNgtkZQM3F/a1Hn
Y5CtNXH8pLAshydh2AUIHf8VgJ1tPUUH1AjwtBNRoUK4if6XyHM3rjOXD3vwCZvA+SRRKCxSFBFN
f36g28UuiaFwiVFECpJBLtkJAd1t1kLmFDD4aC4JBiQwaucmgnhpeTUkU99dYXlEZg46atHMRnfW
TGH6k0Dw1/blijLf2tLHsHxW/iPPciEnIpV77KGKXay79pxTM6YwtdlDHI5THgXV1ur1yi6T2BGl
WQfwJ9pORIapMM8BNnCG3brFpIQZevBLFl7+YHUHq2XmNn27jWxMKCDKAFLbE+DTkUJUnBkY1PAt
INKQ4/MEW+RKK6PY+FT08rrXmTS2qzGnOP7CrnLUIL50Qdas8HErUdVU9oFsy+fe5wU4TH562uBt
tu+xl18W5ZmIJwO/LYVIe/QoB0kuADGmPy15yV5w+d+pPcHJKl4KoERK3LySp3q6HwF+teKRr/x2
h4RmQLsm73IknJwr4VctVVPfBZhUPMOO2EGmLWpqTEaGsEzCaGnu5m4at8OFS+6Yun8LsgmlAG/R
sAThm8uGaqaSVbqojzpXljuA0IuWlbD15/ZEjN1b/VSWn9PACVoxy4usmwreErsjJ4J2nwf154ZV
sA7Zj0eXa2+MgBDWIwhy8aAlaKY7r8zzSwWuy+mpmrX2sMvHilCZ7Cfyqe0zg0DsKTERsHkuki7p
DW5xx8+BSO8xb4df9Esz5v0tHJ5JLbc9GL8r3o0zdJ5K81ixMgr8s6XkBmb17qMva/TApdCY26Xm
w3ZSZU3QHbeLM02LWuSief/FBEnkKFW1KlyGLZ9/pduziYHG40O+1RVelTNMLh0l1W6yF3AohZVA
+HzmmmyCzzJNUqrQNBrJsqAfngBwR0EM93ntmZLgWpXT2FufejUFiHjHrS7dWb0mv+ng/VIYAdtI
nxSCdCB8sozEFRP9xKztYjJZUr9lQGk3RqLDtH6oPjQ5ZFy0d7VSdPy980Gi7PclFBJQrJrr+SZr
iBYXvYEsFYFG5Wp1X9zTSFHjv4igLG2KMW6pRToJoH3fZLyaG6rS1XwR3sCtbrt17vyycklaTkbB
/g8q+em1GdKOqbwdrlP1RG69R7S2AStOccTJy7RJFKjqWgC1K1pVDinmgifLf7f06uTSBjVQ2ZRB
wj6UzIlIPKqiBXdad6zpGyAL5pfZWy0xmFDSUjJCtpNinmHRoXOxNBJ2M7npG33bl3TQXpc3Z6Tq
POUhjtfPmVjvJeirhjxNHhTYsTR0/Dzl4JFNLgbSRg8lMJQkDx87MNkjl/BoMXAotgJ+AfDoPz81
COzXtuX9fsNAfpgBPO2YKAZy1B9KA5nb8rrw8eBcrP9EfIfosvqjtTWXQd4Fzz9wDvdtfLg8pnQ0
FuUJgwkx6Rek36SEn9OD1sXvMSykwlfOLDWrST/XJ/oNZCUf2hPmsEdKSboVwdUfIUKElV21hJa+
Z3rVO9dz03PP47KSM5E//BWTyZqaewHp0FVGiKxdEJvaHACcL+dmH74hjHBjXDzHIvJdVaWob6I/
3XXcMI+/LuBys9RayrCYKVdqIwJtgjr3o7cHoqOoDyTmf+VBELwlMEpM/9mqSIiHXn5iMWaLtQl5
qZdlWhiSPI/lq9a0+SPdVaxEVs/ZYl4GkguRr+/nxVyXaxbVQ4JLPWyDjTC6qfBtviCRK5bWm9S0
gHpPdiDk8ODmgk/FrrWy8sCfnEcUBmLeVJffLvy0edEfMZz/j9CfdpZtGn6SzuQY7kh6qapOd37C
TkRDlkiv73249uxf7O+fPDSDbGpxzmuq4QLPoJ2lpa+cYgKAvSIPTdalBpnHabOnKDlj+2CM95Bd
L1SEQIJQRB8FjJhFsc6Wnbi9cARDhzuu1N9h1b9M+aS0SeZF4cq85JHFWgbDzuGtQaX0PMOw7DJT
D8brJLccXmLhtEgUZDnbHSOpQeCjmo/IUhZ/WPALW+agkIZqFA9MW1bK07ehTA4096rBKSSmOzl2
sxCb8OT98LPLVgwxtfT3BH6GVWI+RX/CYd45O5rFCid1nb3R72QTTE3i/Z2Z+rbGdE21mVTF5Mw4
HK1rWbex9u83nkw1OHX35gXkZ8DCQoDJYW1bk9nFhNtR37bABaGudui2SQqaUBWSJLC3OCk4YVdy
aDq1uG2HFpRDzOtWik+fgGPMpZP4Mn3mjTToO/h1iNn+Kns69PZ3r60A6iIDJ/yykdW1lN18e4HE
dtwVvhzc6eJWa+RNY/bIcQqpxbo4bFWysNp1T1LvbLVdWtkiCrmKubJt/9JXBGQhUGwtSusyNylK
cSSNkCtGwy0pMvKV8R0anXk0JGjCdx7/rlS9g85B9fh3mAlfzT/vRNHgRyOZmhxHZdnZU4PcClXN
dTx77X2Fp5H9xzl6CsLM1Nb2Z6Ds2aWTimy1l1x2zGls/C8g26v2pOonnFIm0eRcHQjJ3M8pJVcq
/1v3FNoMCLpdmXgnoPccZl5kEpQcYUO5cVa/x1ifUVMJU7105Z5iFVWKmBDshZgSQx0oGwbkbfcB
/J2ZjuefhUSK2gZw1LmNnhwSsTgN5DyrUV68o3om9MNPbvKjJzZA91ZjBmJpCCTVzRtOrIBMkfPy
iUG2G/ZwXm2jrA5755XROtfta+LtfWeDbyxzFWBWRH3LEUYsT4PnjvQieQjhZxP9bQZ1rte0KxJF
+ViNqwwji1CZXNI51R+j+ueX2JLQcA2Iz6KGAD0APjUu3hbMljkJ1k/UdArKTMpiyqN55VLq3zRL
juWYp1cFHK2sPSVM+jMSeao3TcophgCIRpfk3849Cn9k3lwduCnryA6dzw4L8x81IcWPTs6OCJWP
+4/koeE+3InM8lHjizmyapydqDpACRDt4mbPcixZoEatygx+Pzby8fVmhe27ycwuodzg5KeuWSwX
wXOvCALeTJms8VLex1ZWyuLiF37q9BnhLsl3YqLGwAXV5po7FLhrYp9ph7sZbYvNz1+RbF0Qkotb
coxqKbm06weHE277ONUB2Au2BNTMwtzJrHBLUZNp9IVUGXuqcnNnOUgThb/HHLRX7MBOBxCZaqr+
Ed3vs0WzSOdZYFTw7/IN0ZpsVRoSNvNlk/wtskHkPH8eG91O6XmcrmnJZQF+wcdNcdQe6AAwbB4N
M2yerBJx7MWNEL4qIxZfSMZe5DBaruY13KGOgoyJEZ+9jCwUtFwMwQQASHnE3qvrJgiToDSdyz0C
zt4RYEQwPao0VNEUHd95c3Nx/ojSj16dxOtYBgqOrYFahbZJC7VxcQ9CaXYe0V/P9WoYq35NaFvC
wGhOofmWCRQ7RurvHoHUqJwLfR3avw5WwaTvtF5f7Lr9wJ0k9o1/wIvrQT2NbDHBMGmSSmMPbJig
VtciXsfkNOZKZtrtzC+lNC/7B+sVogsiesNZ72tezh/voYemRjdUnVJU+nvkhtmDRFAJE04idm42
c2N/eTHp7vi7V6LuGCvdQI+0X3MjNR2A7O1hsIWMPKN8tWNOXB1ai/xmyZTpdUeUjQ4wA//qEwIe
sq0mSzpSc0Q9ZK8Ktc1kRcOG+2dQ5Hr35QbJ+TNEdHnFSi3QdH99mMoICjlyrdcBX41NmtDo8jxB
I1iHMECNgVaVPXbvXKxvero+bXKeF/O8aAtt9eHcF5mMez+wekih4U7RxHjZsSG5u0wV71gDbbkv
MQoSpaBTsxWh5mZYD6XTsA9nFyz+UWqNjxKDyeioKuN1AQ7bU+0qqrI4zZIyVcmITUvPdDj3le8y
8TH0ZpS9nwv6T9ZfZf3zjTV/tABvCdXRuidFWSTn7cADGDcJDMlKIhfBFAprh8cJaKLTS1/2OXvq
O5yVDY3qXHABkfKeefI2b86DaNYHlsRtdRjvuVtKYsvv8JcRWC7OlmO6joiCruHS9QOUUBmLDjnD
wF0Dqh1ScX1BrtzIokX83q+JOo5t7XSGJvsuvGGhruznJPt/dX/GoLy4nEnWEcFOQorzTi3q+P6W
phXTJf2p02JwES4/tbCfkJSqqZDi90wifqMYkib8l0nUxLTFKsW+ZDRom5Y8VJUZdmwd4HujKf5j
TeuQFGV4ttpMbPjqFVewhnJ0k3bsIDsd+el8X3X1EfobCf9rOhOClFBFDU5q1yOR9iWDJGJLjTiY
NC8X0SUqHu36gOtXGJ6CMx0u2UdQdj58LKTytyXffORQ9To6w1TsocJ8ixynUEUGRzhZySOHdUV8
qXbLY3MJm6DhlKjaYWauJKkWPtnn2JeGZJcKxgSN1/TZmeS5VjYwoxEIlzA/VTXjwd0lD0vaVRjG
W8JR0ICBQjp7S0h4+nklqm49Iwu0dzG9Slb0y7lJh1EjEO33wBECVhMUupQBqoLWvzMpPCVPYNRR
e51vvNiEb/Zb0dqpyPT2dkySZqtzowBI82QtsIMj0r/gOlSapFiZfHvBtECcO1ahvf2xaKp4e+p1
aa44BY0ZWThQZCJdV5Jdhz747gE3TSKMlKSpgP9NuB2azzKS+6Ln39eWaJwEua+QE5Jtz02kKaYh
WliUucloYEIqP7LcguIayhBW95x4rzZI7Ut2dFBysyyPv/SkMQYoLqwncoH8+3Tu1C2k2MEsDxZV
XYucqKdBXK+ELQOFyl+PD/fx7rmr/b7jYRdfRMGZNLQpOqMeSnjn94+r3dSK49zCm1e63qcPS3Ed
BUw+rbie0ld/QJ0m34f6CiRVLmKWmOhLr3O8PH05694F63a255Qu+JXyjw3vXT8omkK0DdLiWFuc
Hl3HzLIxAUZy86jFStPg1B5A9lnnDs9wzgy3LOgldUROUNCyhcRpPZzkGl+dmIrVrcjEVwDwksS9
C9Y8QTlsjl+DouStvG/NuThASwE/8S2An6W5bjKZN10zoUmp2ZL4qB7m09ChxqiPcfyjQjultsS0
fsCFGxlMHGHG4aFMech2rIk9ye/KoUDiSKDQbN0DBo2muWxU/o8ZqsWrB2PDJ4fQ3pFm5aPBIaKs
zmqmlkz43YtZzmmGhk6IAAdyOHh6oezAZbmgJm0V+4Ftlq9GZ1IJCT6qbxkWafsROfK42jN0SQhf
XghoeWkqu+hjJfkVmMQ1qz9x/EfDBgPKdwtX6H+A3L8P+RXUfMqF5073S4JyOBCumN7NU1cBZnvu
fDPQhTD/aLymp5KkiAEu07Vq1vlLA1mV+ApzLUtUiHFmhgf6QSyVnJLaTDqpltrPFLIhk5rDx9nm
bfpdyRGtuyt4xXyY9MnOTUN9NU5j/HZeFoIIobZAx9O2nzq+Rq8J2iozh0rpFkRgNJR5hBct8I88
ldhiBhux/AsWoxg3ylXb5/UN9oQcG1arNlhiqmeIdm3rVZrfxks3lxqADWYYsYUzKZ6OQx7YvjNc
0FL+L2vkP/0Fn/UvUBrdqLkiGDTWJLs2iCSqVYvpEqGxITn5hmnMxDsRHf0j8Q5R4zH9um+Z4TVS
7bJAnQ5HDRf+jrOz3wCpZ9tNvC2Ql6WVDHq1LvxMy8ce407iv6lVnYWIYRLrn0O8GUQc7dZt7AsX
Li0dKf3KvVPLkqV+eJ0er1RoNVcxKAAS1OEGB4Lr04WQuFcGbpujntwesJdmG3YTzfXhIA/qIvkj
0/w6LIKme+F/UQX+REo4n6PyhCEdoja+XaRwU4tpwOj/iil21cbP2OTJVXqUDzlTDi7bCqRHrgfN
8gAho9Cmb9xVAFF3iKQatXvS35Cl0YVvJw25Npe8F8Fo3Fq3nqMo65/MdBvEkP37K7agmASkGHbi
nC2MmK8yffymcQKAJKpH56MjrkeoLLUWkx9t/iT852zaOt3e6/VcYt/sWCbkxV67YgbZANzVr4/9
IPMmda2MFRVSgijvO1i/ad0jG/HOPwwWu+Zz6k/rLLdku7GsFZWwM+eqOUeVGth7HwqkZ8x6Nhwg
3zkOY9Sxeb/VVJHjfAn2Bfv9rHRQwWw2I21vDui7FRhtWoWjWAQkr9kMku4kMhm4M0J0TP/G5kZL
ZCVaWiC2yBVWflnPQpLu5dgP+6BhQQ2cWIjkREkCtfN4iniVj/XC2q1QoqoB+n+9CbrVgRQ6o/xU
QvNVgp/hQMRC1wT6Qwq0IXxQxr1QyOXBvBDCg9i7c2amuO0FIWjjpl9G2SFFK8UIWQMcEBtlh2m3
pBBMLpvk0te0wMG8/EVRQpaWunvAZQIREu2ELeoYjm7hrKmVH4e9GuApMZNQzYEQAL1mlH+wiejE
4ikGhl9SnGkmUVmZSy5Tql8u+lgv941pVksJpmVViev5v3/kHhLJKkfR2JCqe+AjqDFuT1Qh4910
Sc+xjEiSermVBamymxdKOGAWwo70Mj2YU5m2vtn6oLWgRxjxGeJYzNB8NisOOBiSh4kADainet7y
Yl6Bs4f3IMZg6XllkM54PuRK5EVSsvQ+Zg5kK3EBg63qUlqxIRnoNPNItIC3I00KaCTfDJvYZXX4
8XPuZlhMWsMQ84Be+Hvi5KwfatoESMdwBw2PbYC9nnLA3LxfhNbIU8wcksJfXKW35pwsQ1qLP0Kl
im//iBrHC0YBaa4hu9aiu728zYuFF6MTM6BCdzP0EZGi/2DCNUgSibz1DEUxJL3huJaJ0vtZemA3
qSq43tplqSnkGkxQ5B3uKgY+/6ljpCcBU6iLXgSzXsJxrD4LGbDLfRbLegOQ/dKUw6xkK8CEt1Ql
3qQqpVxxwUBfHF6f69YpUuWZ0TKv8+XlFpKzW9EoWLwe55UjJa1NlkZfX5hAeP6i73bFI6tUeFku
IKj7lLeTIPOAFeP1TbHCcPFdFLKl0rVeeoTK//NIMwo8vTQYzCoCRq8lWTh4LEloNeJ+2Fheavr5
7IFIP1BvOZe+lxOJQ2k+jEyxim00AuFvc/HPcnO35hfTeuE5GZ8I2NV5q2sPLJrs6ESwUR042O4k
baPOvOfVkD6VsdIxIZEMgJpSpCitI+C0tINXTsBaThJxsTHCrhEADiEx+uLOi0vNPJ0FNcMW33zs
LfwQWZZyTBLITIFDLcNnlk2VnDZAkFYuhkP++yuMjo14Xro9HZEpmgZhZwYpNuqlOM9y4OsuWCxM
V4m3zv6m3KMT9waUtd5pqrMl0klfOPyOgLnglXwCw8rBu4Zu155VWt/obGSi+2Fe4G8UOs9F2Nr1
n5UiJn87K5hrtT4bbhnC3jYJc/9rrdCnmumU3Yv+tP4763oy4evXopQv/K2euc7peKGpkntvEic1
nvlkm+n6UOSC0IxgQ6zi/HBk4+qxhT26cGSqLmnvLrOobG0CWfTRjD/vFvpUo4dnKaWms3tnZksf
/+nxcyDX4XlfyKFUKS3vnTlWigP+4tsqiRmmP+t2XlSMLAt5hJS9DQX3rIYKhxBVfGTzZqYDLAEH
r757R9w2Nph9QLb28xnDU6rTc8ajmMfGQgcZX+6fGTCACGU/Uhlzq4uTP0zhviuv9SXzN2yzvlGd
pqgu38ptsAWMiI5G6zQDayRgquCrYgfFZY9uhFD1KTjHwQLApq2OBrhSAZ+dPufIJVtnze1BN/XJ
7oNQxFUmXdNa5ICGWvs9jhge3tBZoAHq5hmMp1uSbG+XXnoH5bedXj0GJy21c+jHyaxJgn3lkSep
WibFOeC7moCBxMjqTx+j4oUYRrI+mQ4rgo/8zHz0mBX9jCAzLoV7wzOXCcdrxC+sexSPz9E+CiAk
7ScXcffX8vTVqQn5DDl1RGMBfLELOyDJD0eQ9qCgHLONmAMiUMmmWluG/zIGJKlfiZpabFp5WKc8
ezreGq0aNs+i3n6Mr3m8M8YTEXxrfG6Kd/AaRUN3Zl+8i6y2zMCcWQIAhIviFfkmST46tllrMLNg
BUov0UT8iCoEIm3QsCXAO7AdL1FUNi4nOsE5pokU8vcmqvfrs14XF2SVCbuSrJ/Q2jfBtbRxuRdN
xpOVixpxNQqL5cK+ViqlLoPLHT5LnNVzHXeEV+y6t506AgXWerJexK3O7pWzoFqUBhfeMsQf8AY6
xTjpVIY+2pM1WvZxSO78/eJVqGkfsfFB16Fjb60BMz4h+tYgEVcW6y1BfrE/7z5iPwK6nqFF3dLb
wdjDTrXhgvbaiqHrLIWmDtflYrwL7199sz7Hy/OIe63Ng5wdb/Yeh8QFhCsUceF5Y0+311OKL1OB
xpYnUr2UIEM9Ag873AnLEEM1e0vH0mTSAmWraQHHJu7V7KvNeQtioUzlg+ADsB0zDY7Mvxbz2OdT
ywliycsZmY1TdHAHhbBpc29jBXbJeiTfNAh4TacrrJ3WnS1+8g83DtET9kBugD0rTRpi9ZElto7w
ie8jAEnx+h/w0TGDeGRZ9E7/PAAFgFE34xdMnquHcqnRHc7FBQfKxX6UfvN7bY/oqtTZtChLp0Z8
DlCBV+KHwkRWEvaT0ztpzSrHmxuuEoa0szqUp7yREx7E/eprjc0X/EixNZgWdkKWjuADDbScMUCC
CLKfkP+ESVlQF/q0Hzs5FdlzkmWBh7r1gOlGvQ+gzQdTQ85ZX83kb/kMTX0gYsqLV7EN7h9fXxyM
LySCv2FJdK31cEynUJb+EzNBhVvZYg1ConFXIb+fWYhFCzzNQguwn1yezOTFMH/WSRNQGVTbscUO
q8tOoQCmFXG3Lu7j8KLNZlPLiBhvDJaWPHy0yRSEFNmleWyp6wqhaYLW10VoJVBmWbVfeU+3lh1N
JRmrEoyprVRhBSO9dqHt5k/1UV8UpdcFZgtY/yF8NAHQRPcuRHjPnH4yilSv6+ApMsmIg3/hitiL
2eMmd0R3gSJXfQgLzTX7acx+KcOHQWI1kr0Lhpes1MZ1UVgXfHHpJr/Dal3G2B7znN70neEaYSEy
13nxSLFoGZNhxjQM3kSuoCbZ9OTjnWPyVujlBNHirY9dgwJ4980CmUJb3IQs3UHl10DH0I+SydLM
bqlhvjv3VraPTl9e0BsQlT2kz3jGtLUBao+L7jr2Qbq1fWp/MNqXU1iTrz3PKv4O3euoR2hYmZP3
AXsBCLZtpkr0nX5zYaj5pjl7g+x4sYvrfuIb/V9AAfGMuyOmuYNv+Gkko/BDDme81qdwc8JhxTTz
ha9SdHTQq9hynYP4cyqd5/rlLzM7LJzoUCbbS1uFQZRMW4jT+raFznUzpFxwbdi1NbHHyAtK9Vn4
HwJ7sCFx7v5KpRFrQD4lQ7e9XbkUxZP9R5p3C28OM3x/PXKwPtj2GBANOMrtPZpbzDDgj+Bjfk4/
meQqH488ZlPs6Ey8c9Y2Ug5Q2BBsAmEbsm4W7TmV9Y2Rz1qnGFRU2O1aAhI7jEGPtQYQaiJbfShy
xngcgvYt4ZmvktV+3TwhI4MC/44XFmZ0+9SWb0QIL0pCVj2wLo3mhJOM0u/hsxopVE+S2kBEzh6F
TUTRIX6xnvz858oeuDxAEaAyhKPAl6Rqc9QhZXS9AdKqQMkzJ8UcM6MR0bkTkHDlhZ1DWXtROgxd
mLH6Tk4kmwu8wOYJJPOXdD8tfL8teH2tOcHWQlvUpGHtzZKK1QGegAtTdl0+9iwaArGTtS3f/slN
NGzqNg3OGO69Sod2/2NTP+PRWvMc+3RM14qLrwPvbfxQZbrrJLgm8syNd9ihgFj681f8UzbnTFiJ
4U69qkLGM9LKStuPzuvT8EM4DWLZYUI/OLF6yTm2OLbJBX7JXPA2PBpJvVjkkWzC5z+Vc+SPfBN/
217INnlZYLxVP62anssUxXwl6dtHNY96hky+oZTz68f3rRmAE+InNkz7FOCn4sQxpE2XTRrR1Kwv
iRVrK/dys1/IeWnXhNBePJ3xXd/toMDSKnAmDSChZwWOt8WvQdk7F3AbPjMKi1d1aCtbT9ApO7lH
FulaHCLiPmUwx+E2OZwuthM10BmgIchA3P8joyQQzWzAwNf3kKB9M5/vRbRgI5T5i9WBN83YuYRD
QzQWioAo9O1jdsJde/rtOZ2EiCkAzKTix22cZW6blYwAHfVVvbuiFQ3fSE19L95yAZ8IeA8kw2qG
rSCJUnwtxTDZS/a6wdjcO1chg4EjAeQ8NvKY5/LbAlghme22F66xHLMSQkHtY/J8UsDGyDhu6dPf
k4bVGi0pMz5krakUyHVOJTBLAkclQXba29QZvpMVM7W/yP4hyTiiLXZc00ymzsN3O3ac9Knwwt1a
ozrT3zduIO4s7C9QY5ZQrnFNH/2jzK3vT+vg0dKfL+xxFkA1LhtnJ/XUKB4F4lJUR0eL0oGS43Of
oC8ZLA4IaP0PJ1rg6LSewR/NBeC3GlDJrwrPI/wv/OMWjSex4kS6OEGSCklX2nih4ksGHpHoIm2x
HsD+RdV+oF8wXiKNDbFrfTZG6WqN2GEyJ5Te0ZXDNOunhd5yiA1mzXhGEicXRNdQXublUxwGrFHN
kLhCUNHCMnx4LiU3i7k8dBPoiOn9IUzUv1uXNuEdPh2OKPr7zsaPKHxpvBKBObs/JihKlKYV698e
K+0Y7yvjQ3SKIBGTMe1SSU0sA5TPQ7j5AP2tDCcEFHAc8zpeRXsClQS5FjLmEPgj5Vu1ka4Jpk0W
OUlYdSnds7PBprlbFoK9py/nprYfg2BPT7cX+RWfpIapnv3rjQ+hNfG940C4IS8VzjeIwAKVLcMY
bpBrl9MWUc2Ah/KnxEG5AxW2EdKlEgfxGx5N235djuMF5K4f2Kx69fm7feeNaeo/vcnYqvAiE928
p4oT2K6GLCWngdtWIP7DvnTSRRCPK+tgb6NycxiIGAMW4SCwWh2RoH9uFId7eT0xr4YblYB0a8fA
GwRSOQ8PJE2X1TAVXITZe5kyfZ47I2IbuMCiagiGWdULbVZjUeqZANZZJXEnPm4Jnq0PTvPzBqlT
2Gh/KSEk46B+tyePQOa/7E54xTSfBfbHRSXIYAfx3JxoVljzIWtOWMzy9CBWU5CEbnV1Tr6qfnSR
lrUfh22rYPWkf8zcjYxz0XyzTD95uizKu8CEzr/mtjjkZH4ljYkK6Q9zyFDtNqUuafKz+C1vB+in
Gm9mmZHQNiOdUVhQyZwRXyjK7ptY3iwWwrMuBpvgWDmLM2xrLXAtxgFIYzdVrYZQIZBdrOYkJBcf
EwblrGmIgh4+F87tA14mKQSeoQ6GdTEEYlET8l0vfLxu7/mTAaAQgwOsXQpSpOrUv+Cve5F8KrUf
4tyXxUMb3itddB/qAtSlshP005cauzVBR1Kl5PQ0FwvfwvOja0hXs9jurCsne7emdei7q9PBXVBH
QGkTaXtMaD9MqC4ChKEWgRWTYS5Gz6nOwJ1ZxGvxeWSYuIGU1eV7hS7yfIimhAACDQssHjWXoXmw
+rh/W9Zug/j6MmgkqH/n9qQvelHwUW0J6nevSVR+cXDsk7qNvKZiVB57sqCSI4Uqx5TJMUYG6CTT
zTUqxKGArQAhfAzbOAAdKk/hACfyXAL+/5whsk/iIrCZgFPe+tFtl1bJE8LXzbX4SSYeHwD2iE1J
UJXBnha8TDOTbQp9ptg1zfQa8cflNpty2TPckSJzYneM8uskPWvDiLIzyxi4/3Tn62s1/Bdasa6Q
DHFz2QNcrXvY2X/ONVazHj48QIxIxSkuZszKKG5VMUEmFox/3uUPRtSx9Zv0L8RpzShdpfXejroQ
9BKZ5u20e6cyDUmIV56Cw1zEt+ijEaLwg5wEQwFpCT6cxGbGdCmBXHUyzfUjBUB2j0MG488NwiZj
W7ZaQAxyJV4iCR6J4quJy/MjWJDAArMhx9vvt1499mjRVyoTGFWRsu1Ahc/iovN8xHo9UBn2zZuZ
Rae8Rrqki7ffIZ14c0eOUe/mooWIOFS/JVrE9sJSls2ORMkTLvb9a+tRxTYonvm0dxlC14UxCdK8
5E4LUn26tV3IGpTOG8dWj3+5rrIxhShKrJeyaFVkJ8HqUzP5BdrFxKL6iTBEzoeDjASrAinj4DNf
C8j/tn3/xXLXxGamk+zADzsE/LMi2zxM02xYl9KFlZVT2TRxK78Bhwr7M3QWvDzv+tIlUtaYemq0
s9Ad1wW8r8zSgPFT59viyo2BLIHM4uBdIfS/CcfXMQnhv47ZBcOeQiJcigL9KIOxt98SVFYqKne6
5vBumSYov9wFRZ1uXws4g+NlSnIwliYyiK4WLhPn3OgVsA8/TrnyBJ8W9picxYFihfrag3MKTSmA
tTIRNKIkCh4DgSntJtlBuvDRldAZl45kyKmFAFN/aidPVjXY/lciEgI2QQnhgAQZwDssXTZUJ1c9
IGV6A6I4V9X0rcqNumeYllrNpgCLHfvGgCWWxqQK4VM66tekL7r9OtzS0kRZCabQ+goZWLKRWFce
9K0OrT7m3xk6qYH5g6WVeO4/zW5YxhNb1TohXoEbFHCn1ZtZ0I9xph44OzhH8QrgE6iF6aUA4+es
f6pfs5GLIqtvce/87//Mg+tFYQoWNBVmbjLcZ0J6L00ghRGkg3CSNgbxjomFTC7VQiZVPn1Xc5z4
drnwIR5/LoQM4FyfwMx/+A26eVVfPvC2jHGV//2umcV4KMiLl88s/FCEYHWQMIf7AKHfd6bXVgxE
q13Xf8ODjEBguUKINObObAEHDAuEk+9zjs6MMbFzJcj1CGeacxpJVhVQFhtM/fxMjsMmfgYrBjki
98wkmHRE4FkPUI6KfIUqc+fBiXLbtNDWzKfzj625mUpF0ZaxKs4Eitb/WKL2tIj8ldYtJt1C5z/1
djBj5ZMiH9vxDK+43ezKLKG6A5P+eMXGIoHNuRVYQdpac19j7Y0S6fV465awOU5ZmEN+ewszCyhQ
lLhW1akO0qOswB/RoY4VoUBtzKGcHlKPz0Wq302qdJZ56t+3dSisxPktaM/ZhvLvuX39KXwLcsaS
Zw/72sGAMwUYsfsCc1jRK8KUhKMsYpUmTic6D6mkdR9fdAc/Wz7W4nCYwSzY84HxPPNpO/8qhYbA
aBfTCqwZRaO9HZuXs2TMHf4DuOJrqYACERbmKxNtCJ+H8THc1zxV8o7OVvkdlhUj41jWmw7oJfHJ
69aOIwew/SLS0a3qBnmoB3xXbXFm5usojxf5NUn65YN8XbO1JGjiNDtcZ7hsUzQqljBCfkSBKEqv
S0gwnyVjhp/byKvchNG7g9nJ12M0tzaxrr9KV5rfinkaxGfF2zkz+heIZExuKBvhkENITFnXXJua
TWkirZ4nGQKtz6E9hrIJrgh72vWwNMJ4UkJRylkfn/1woo6dk8/irPlitZwZumuncArKAqd4fpbJ
YvHZltEhAtinwxY0nzl6ZkEHs77RYjaZHH3qCcYdZdZHoGIwfkOguYYP4ap7NdwuOO0uFtpUzhMA
QiRwgnkwSgKy4qV2k4/ybwiUzJLBS6vTNLZBbVvnAtRK0BVo1OqGOZ+uY3unGwb792OtUVQJhpoB
DeuGo1t9gRgf6vX8zNHrOpkcI9m/s3fYtaoa6FQ1oaWZ3b2V1Nmczm1ncnH7PBQVWkgNNQpcpuEp
LKgv82gMDH5QpJPuMLkomMBuqGaKKEM6yBA1CxV+Xo9XQD16Mxli+vZo6JcGholD0SahWudL52gd
YiE2hKrdQfr+vvA1B8zSNpr8rC+Tpbyk2ABL5sArObXDCVHqnhz8z7YJBYsmV0hEwLJiYpti5K1c
OCMGA3VDZkGANqTFil8bLRNCawH5KcO95jkiEhFPl+WnghDECmEOSrbFN2RWPUIzA+2DEHenxQq1
4A/BNwRLz2LxYOyPKGxcQEQt4HRYw9+wr0C7fipKUicibeYQSBqaLNqxsNtGBUQ1KsbNTLrdQidQ
qvepGRTqZCcXVq5FSeZ4Z5yE0gEwSSQVhS+eEqeXbhmZgukeblZBCMs1FrDfgXAP5wRDwktLYY7l
Jw8bQN3i0WtLVXjvMrPpB5MQK8CmnCFajrJK9MmExDd+5jImQfbB2RuhnY3861oH5bEa8MsK3y5A
9ZUv73dhEwgbKvts1qAlpyXTUI8CT5NUo9aTGLF8DbkxDtZ4+70orLmmJMkSJt3znk2u6SVwlqmW
aqDqdNocF/iTgUnD2PnhiFqwIqCuTKC0Wpub8OHd/ZIhm5yMrNwoG6tHJEIDMe2Xpz0L5b4RX2Dx
Tv/ev/6oC9eUTY7DUjN37FL5lNfrVFZndBwSDte6T7mSSL5DE7AAahfq61BI6dFFeuV4xtb39iMO
52g+GEwYPDS0Vse2wAG3d7Ox6XG3T0JAbawy+k1U89aKM+8EXnUAeSgdJFhu/buo5Eamp0zBydy5
Zy/28bs24CPC3epG9kNYHg0RRoVqlCKyUCXEAkAOFnq9dw/A553jFTtrtVNeXzCfv1RjZOrpnAnV
+s0Gl66MX6+5DeBDm6t6ywOiITqcxV43GPL8ILLvDDonVHA+HDD3zT13lW+fM815gNRqf6bVu1Sn
agZ1Fc9o8oMENK6WEy9TEOBoslnrRtVcub1KkHttA5TeqX/7lylkJmOtpOSehXADRR7aLbmsaQEe
1zpC6ryJRuXb4BmLrhTjy1wIEv6Fhf5ET+cQN32ZT6P0XElTVZyZBlACeBx1/lVY5WAjzfML3sdR
4jM0bIbCMPb/n/xuO5OAvxTcu3TswNEkK7exzhf8k1P2RcQ1IKpWccE2tnZNUvHAM04pQEfO+Qfn
2cESgdfn0yDUxxKm53Ttacn288Xpw86UCeKMU4pNt3aJ7epz5rgqLr25XVXuVpA3CHVyg2FnwNyM
k4eP6IcJxVR55yYqConnr+axJqcM/r0s/20nlnne8ncj3QbpfBHH0mTGOncspENnuh9ElM+jRfkX
lemEY55FwkHsYtP2XalWhhN8ZqEVN9Lt+WbhzNetw/D6D5HL9vKu30wECDQay13Y8Xb6jTYUAf1U
r1o5BzvT4FlRTtupDRZaifnj+3dGbNtjlJKx7TxZerDBZVl6yt0VIWgGKtFbTwk1Vub92OrS7lRE
+drVEK3FxyW+8n6NBfqZ/DzxYS28zA6AgXnE1m3+p4z8yEMooa+VE/2QBhWf3cKT332YGfH5eXjY
VWBo/uF3yXteJgyUyJM7NqP9fCijDuPz48tNgVqfh2cpUczhIqLJl5DVkOKpSclvggAQ6MzP6y+X
Rttmpp1YLfTYnttKwgnh5POmNl8/Dh5ky3sPicaCpCts/3GpW+PvxoEW8BTsjBEwWaKXHeT3VGAv
83LpA5NpwV2mqM5mzneQkVmcWXiakIn+I8qwu0XUjAlh2rMY+xvSUwTMjvemHFkHCxJRfEo6YILh
ngjhhhhfm9thgygx1LMcUH4E2oQa8HlLt7tPuKCgBr+BS+tKrXN2ONJmo8uauT/p9qXa8YXj3ncR
V8QRzrpOEuxWpFX83GJMORxZQbPXCYZpUO+e/2jjxM8hdJ437HQQXOABZ6FhzZLrJ/7ocvbt3Qdg
OE5FzeqpHIb3PzIbc1QQsTs5Fb6D0KCI9GllxArP/Q/mU5rioKn5vGisNHLCObY5MAPrTzFsfpdz
ecg1SslZHAzodYPXYjcuzPz6ZgNzZ1OfMZ8f3mMmqGP9hKfMYHDiGtFgmfzr3omIPlc9O6XDU76s
V7xxFzrsL5+JlBZo8Bfn1JB60RDAaB6c/JsQ9nyLaY4lyDVqHwpr5JvRrt1xkJbPUJz+s+O2Gpct
iVwUYaZErq6L4A4nZEfTnKunFmxbUq7ssHIn0rPGnUDHCcfv3HcO7VqSso/8s93vQYJf2f1UZJPq
CqZbH8VKjsufPgoxKrTtlhjjZKLpfCxTd8VQ0AivY0PjDI24EBlS4++2mXia7s6Pl/zjxSbBSDsy
IQE8V+lVfKYiW6JdCTslNP+JC/TYCyDRMlCiGwLUZv72lwnbokNWQtovciKfaueK3O8xLWdUqyCC
5MV3b62CpCAYUtZyqSE7CAYSg7tx/jcDDXp80maoOqub75QgAugiiLjl3+HMHNIkKQzOZFJo00Pm
nOgMcqEx1WCifXxiSpDrrMEeqMwmG0hKYWef8u3D5oHMmrk07pLaJJ3AE08+BE+JyYw27+oAG8NU
6SBNHPtkY9KO/1uVPRIdlajdDngAg3evTPGhJXxrUuClk67eDF08DNaWZd82kII+txFhV6g2o5OV
izJd3mREJNjehKHgKIm1noYEWg74zeZPVipAgVCL77sMsvsOn1SELMBQet+GXdsd46NezGWZen5t
UhEX3ORIhcpEFcFxGx8MPh1hFTq3dlojsPTZ4zQ0D47st1BB/GWGjmGOr1lFQAmC7NxQl5LDhFkk
pEc1oFoDYQ7DG03H9vzSZ1FTWtdktE8FFuZrH1ynhjBUOHBuQTUJelHPDQ6a3rroNQzk3ErkXJou
8arhDMN9Z53LMzPnuqwWO09ty2t1SjV0bWoy3DLJycHCbnLPb5RzXx4WWGBfLmidB1cqS/EuBrDD
6KfHuxt/1hUjf6LzJtoXerhhf1vXJdaZR1Ta3qNu9LpjnOuoBbo8odUD9Fv1+32JTk4CjpPoL77i
1koStcSbZYIfpBpN64bo8lZx2bmS9B97qOnb6g1pRbfA53eXzdtVqi4z5T58IGJkMhrbUYIrLF7Q
krrmTuZmSQEOfjvb5819+yUuJ4eNSqcqc8s6LeK/RiubHxNFVwloTq7ZzvnBJ3RYaPhjvAA67QIq
mFeGDnLajjkZiqNaQGmMbVPKKmwU8TI2a7583qI0qwFl7YGsrEwXNJx0Jf+VpD8gd63+NW/+ZpzT
hXVv9NuH4hyGa/f2JwFsF+Md+agMcbtcQfBQvKb3OcH+CGCa2OVDEJvysgpGC4c1jfMki472RWev
gdXhEUCYQCPSPwYhO8KtkV3V0+gxxDmogAuzkh9ej41RHaL0wnVIkDldGwGm1bskK3gSC1plpp0V
iZnGAho3WlOa/j7EkhWb7LGTqBxcXjNqGqFaLbNMKlEQZFuMnaPIbhSQQVC/cpQjVef9YqD/qk+N
W0X1vWpjnwy+xA0QVLutDRNN8vozf1iX8clm093pRouPbDjzp+HsloKjYIfJcwsylM87TfjvQ8u+
sxhdYekyniLBLzT2RT4iHtkyrY+WCFIrYk+L+cGGCpTSanNOUurNSutlqTtd6A6wLmJxmO3JvAF0
kd4tiwOXDwn8yfJTq4XI0URGo2BhK1cleVOJI1992SeAJJ+faDxkZmbuyossR/D5IUpmNAkWeeMA
WOsH7ayJREKfZMAqxepUaKwm0bQ2ngVXXDW0Typ9OAKqqN+wcD6+wK5+3EuFHefBxBODpWUxN8HH
srIuD8VQegfAkr2mKu5mBX8w+3qOejg1//dNyVLo5bXrdESEWkbZ4OXdUCQkpXM4O5TwFkOb2dnh
43zEqC8UzG2lAsNXzFSeI3Gk7KNqlbvQE4qFe/Fn8BCTgx+1BV7ezLheleOX+drtHJJ2SWf54hNC
JQTqTRrZUy52DMeeaAIfV+gjKyQz1oWHL1t42EUByirot5CwIWO7X3mNob3YhMZXzeV14gNosWQg
XnIyDVLV2h7KDG1cJ5OA4t6/LYaGXo0txsC05EisM74h2EVpGZ0uIzPRvH+HeN6qrcQuJeShB86g
uW5a5Inw1q4SK4MtKkJuXKyTgCyj4rNnLmVT8Cnndxw6nnOA0h0E5L+FWb0gctP1EeYRuaFBj6+W
lEofuLjDUUpnm5aaNjXXKdCy82gabpvdrrTvH4MjB+ScG8/GadT5VP+KMfcF9QaRx6H8jnRzRsO1
e0JzmEgX93f60o80LqLva9He4esPMX2wwfBj8iBxqDnK7JTUMvX6AK56SgOlS40ZPD8hhB3n+//8
aROPA5Q0O6GthtsyohiJKRSu6UmK5CdJEd/7jO9RPUA6OtmTTOi3tnDKGw2YVm/xv8LG1zLkXNDG
2v9PmGHD7kSdXrq46W48jhOfyzjgMqqdUyz9/YSHNMR4He2zcH7xX3Dnouy6RvmAfabBS43aGa1R
4kL+vZDR69+OpoAbtS6f9WfoNS+y5kqulH6OHgOSAsbPEBP5cfpNdwXzugEg3dAbyqTYW1NS6YKS
LAwQa8QG+ptNLixG5bGjF3p1+fr7XoO2qqpySSEyYxVVImkqIJMIhtfY2FJuZU/871vRdAAnScuv
qCw1QWJnWBbeCzRoyIScUkb/Gy+3uMAdtAnd2XGdDttLH4R6utDSpT3CrClMm8K3TA33mgSAXOby
lVAPJpEZ/S2oAULJzvIqu3kMnfQeDtxBFaFdmYye2xCtwtXVjFdiDgkjH39qkZrjJlKPH/6Te/30
cYo1ciNgYzt6XIfjFMH37nGFnj2jxMogbBYguFPFlzaipav1ypaKG4CTjnlKexdrxcWoT0uGwAFt
zmSNb3lrUlSTrw5Rg/7ixUfC12WFh9nFp254LaN1o9ipCigTKVnj635eYgLIZCkt+vQHf3Gy1Jju
hjyFi1olPLNk+nbRPePQRyhYGWKPxblmIQilC9AA6JBTGP0z10Atd4HEDDt88hqT4igkymV/sq/E
ZOi6beFtDeZycOt8sOfcR3TRA43djNGY/wRr50MT2TzKaFKwzli+OxtSUenJ6Y5mnOr1d/evFLVs
fU34zgCFrnMAgL/xmnnFHv0CI9D/sczabR0sn3+MPv35/mQa1wFJFz5/0kDqIk2AseHGH+FZGbX8
O4weL+5IdfS+fPX9OZgsP4ZkejZp0bDb+6Veb7MjrjTy8951IjLjYwLEP5XzCa0KnATYIIt71Z3X
yXQRS8oLZAIGFhaxbqnnh8GYXVJObFv+UIP1ZOl50ldoXqSSWFseaitjxbfUidm/JxdLLAxPM7Zx
E53IxG5pO5QQhcO8RYirCkSx8VXGQsvM3cWg9I1nIk1JW0/0JQ4ioeMG2cW+5g9heO6saeGzADHx
SNNXpyNFxG5MZ+3AR30DSfAgpPfEOjIC0aErmknlNLwADttkWRY2h5AZnZ+zBwe6/vApCK1n6y2+
3IF+UKlbPdDk+su7lDoWZ3JCEWcO9kYXf+Yp8TQe3Ius3/OFH9fDVsTKsQ3C7bMHKAHwAvMog/fW
Q0fVAzAlP5R76r/fnFkxUl9y6lV2KadZEVe8bF8Oj32oCc+T86Vh+uQ0a1uZJxBjosPSV4M2Khgr
izd1Dav8U9cXGzuWY2hFFDGeE16em+5VmX050NKVQWR+mC+5LM0avLczvu0rFAqVkaZ4VZe44MP/
5wGS5zmzZo0Un+XxkROeZEuqtVjrqKckPEpaoia6M10wrUjLA+lRexnQ6V0849Oj9ISugNd/KuY/
c0BHg8i/fLzUe4+wwV0LYli6YV1305XrafS1xOzDkbs56MS2kQ9BrNZshuMyx2ada+VG0SuO58HN
k+/vTSmS7vKO5a3bkw3laXjRZlTmFVQPMNmPzMBVXjwL8Hs5nJaBJ3wIprrwZ09Fb/K9FNBqfuTp
XeUdIzLFI8XEBif75mN4wJ4NjzGzSllKP5htizyggjuCq/wtRvWwd78vwg7B7aPfiM5ISpsr6Kpm
SJV4xqRpz9g7dqSJtqSrxMKJbDG2ppiwoaG+zg3XCNq+k/3Idw8/F7tUdL2NkzokjhGf2mbbV+Ih
alrHCKY3XweRlfRuANMRZlSPk4t4m9Q7mWuRN7DShVJvACkaWmxnR5RAoD+KzSV5KzmL0NIKWj0l
J9IIqY42fshEM7kxANESgsvNMTUPQfBk7S0eDNqA9+WhnhLbfUOdRMY2l0lofUmGdoN1/FFAaf8C
WlX/MZme2U7wsDNnPs9bw5wIpXzP2N0PBJpjfIWnwKQ9hfUI2nOUHDVa9VKv7bf1VL4Eo19s1ige
NIo1kYjtPL6LTdkTqqdAPwpdyFq52QcUHbY91cOCmrhltkypWrIlpWsjAqDEXB2PlZRPAl0IIhGT
B8+H5szmAPi/iGoDoMlJGeVdKwNLMASQgP9XB6mQtrwZ0SuHikz9NPTv0+GEIu43RsMRjXcLuUDg
iFOGFEfdjmsG//gFKRd3r2ZRPFWYHqa/da43LLAdDYnXxSYV0w6sWYbC9qBv64oux4GIZiSPPfqh
CLAJCwZV91DIX8HWAK2YdAJrYegYTFjC4Gb3llqlHKxZpFP6EFM7deuQ7aCs6Jh0dt37SVzDEdF7
vWByFe3wkGUnAkqGLEYWtJyDhseavuzoaKEy/FA2XYRhmYgii26uF+VBuDVycEirYn+5vJRTuSje
RBgQnwZMynDixsE2TLAowVwHwFnzY53Lzfwux4W0zNK2fvgp+eiaWrXKxVs5vYdzvskUdEKtQRM1
OUtNL5n/TdK76qLRngo47yjsFmyMfzwGjwbwNDkaIakyt7UsZi7rZoMFV8dUWCXmx8gS9ITQQ797
IANFClTFdkiviwu71bQ3t5tfvV9/cqhxXgxL4Sua9fB7X36dcZtqaRVdyKevkT9eL36sxC89aKdP
y5pKukebFcNFhAkP+8Dj6pQKBKKjwPXznUm4msg4vv0GOLdXCyortTkNCxu6YIrTZOotEiKA8DuY
rcQlCeKg3LhWwNMmoYWfKlHFFIIQe/LlGziwJFz3slEPKbzeCd139ZV+EkmOKJVWW/wzjmhAGZSR
BzLlKXD6Q60xsi31BJ4gaFPuxRHR5Cpy8hL/zwO8noGhhRqK1StkREvQ4WrDOV28dc6hqBfzdAs+
0Isb13G3VsZW0ICiAmv+68o/MpdykO/rQHGf/sO+YrOyLNrQDTmaoqzBvikhEKT3yILLUY97Fkb4
hKyyVIzL8VwnSklmUoXng6nhUMXU8PSjSODC9SYCHuH5XWBmWNm3oKiWBU6IcFjGAn36a9zpMUDY
jt1GefUUr5L++KqgcDX+P2y5SYg/rLexLWpyLnzVW91BKdmCOR6DKvW6txOhj7sjHah3iJSMKxQw
gh2nH1dUTNiJAjY+3h3p/m3sNMIOrVpmq6VOMI5Vdpb2rBbYGj9GHFqpEvarXGyvYwqOTsbeHhII
S2t/MrohV+z0as9yy80jWvSS3JJyl20EKARfWcpLbC0dU3S5SQlynjTz68ysC5j2FTGL7KgR79zi
zKs+KCzpCQzfym+wYmC8Rlodlhe933HXg2E+dqnUqucICN1VL9OoF+bR8T3mMDyH7L2eRxr9cb44
1BNnm27O2SQsLuLlyc8UTKeJtne+FIDfO86PiRjZ47QRVz7nSPwPFd6lz+eKtM9SOV8D3SmDZY2c
86Feb4D38LD9Cfrfa0IZjiL5SmlaB75rS/gkhc2s/Sbk2Z0nbnTVhrUpGBLXACXvvYP6zUBGnn+i
HdKvtacI5ZYylohc1iGAN1zGIwkesHztQbglSED4Vv/8+BSAIE66lMEdmvIrJpw+7VJB9UslBIs7
fjeqjtlqOe+HQnHRtRyr9ZHqPCqu5FsYBCvTGprrIAxOIMCiFwGoow4D0HFS/fA+XOPDAzf9KsAJ
y7XAea1KsJDpBfPd5RlvvBSbZvGgMm55RILNVx4LTJWgYNwhGPhdXmCKI1H62qnsfqbY1rsfh1vs
41b3y5ZQBbvhzd1lUuO/+eyvbD2zZugS+31DKMGd+w1GdfPpe3Xw6fHLCI8EA0UO3FBtBw8sc+44
vO9Dw4y6eAzt9jZ6eIJbT2BOVlZnC08GVLon3W/8pZQchcaaBU7AgORFktqD4UnajJJiEOw3Zr/T
IKmXmEMMfUg90UBxcFqmuOBhRwz8SklA1vWhCt42EeJWl8B6m+cQWW2NGcy28mXEeGtSH7i2oRix
+FImmmMh1eDDSeihB2WceE461e9pSHwSdJp/B5tSDr5vdAi09LULQL46Im7+4oxA/frSS/Wgyq5K
kQJdOFzKRBOPEgVlQ9RCQBvam3qLwbXoL53DScShUvCeyJD+UsCQ7aB+V1guPqCTcb8oWGS0I9KX
E2TqujV/qvOZxi1qdCCBA4ogRIuNtxWtOB7caDtyQTgfaaAk+Bq1aDj/pj0Z6BnvJZ91Zk/8qBzq
uTbwEXkQ3TDfnFSdfGpraFcD8OI3jt+nDAJxwO1ExWvQW2UHRmpkF9zU4Tc83OF6ViNTG3fnGREs
2Yaljyabcd/CFLrBX1vYqVs+Ea0OfYHloM94fCpPkECvKmXLHx0xDOwexc9CT/5K87tzSASD7oOL
WIhBJWsgly7oH5ykjE7rgkBhM9Ft2cT9/hylK/EBymnDvC4fWSQYy4PXE7JTM3oIXIFUcCQav/C3
EOySJozeWYbVcjZGkPQGN9dhCF7CtHcH6vkBABYzQqAkvtIzcK771GoF2CMeE8zKpRMj+oh2vKtb
Lgn9k+kIcABeMfX+U0cUT/jCtXGt26KEiRV+Gb6vlU2vs+EzJ6bfNHueG2B7p8UokwEk2FskiczH
FTbOM9USdfYkPlkhnxxTIOrZK7TsE5hn903q3KjFbmO/VWPVMxpZNbAHj2TUdK0ynAZRnYgxhfSN
fz4XHn3uxqxo+Dl/+b8FjwR/AcevYSYOI6gloujzbn534XDuOUaBGTgvoGXm2NeYYihnnwBeJYoU
NRBuCVREKVGSsAj/IAdlrStTuqLFnYTQ2YnFC4ElIYmLzSEGEefUwNXR6HhE2sF7lxJRRHpM1f9p
p1CanqhYlwIEFsjLdH6S2ekW/OIPKcXPZxgRVDuA4FhjZongDAWSjrPhDLUAkZMRt5hJOA38lHuv
Jezyevj/xjWBCZd8ncEJlmb7e8M7IEOReqMEG/nWFTGCSFX0POzT+2nBXHhlCJtzyIVi4L9EyKzo
uESccSrwj7YwNT9P1WeK4VZja3S376AxGGPl2euMDXtykceZq8T1lRoEmZBHqTjfcmRG1KxgH8Sa
QQrE0PNi8H0t2JGn3aNpcnU3AEeEcBSlNyK7rOu1p+AmXefGgK+P9MwU6zvaNUOpz07mgUiUxVSI
Uwb7MWBgJnvYxgpPPV5eSAkHBs+IaUGvDbfx+z73bgx0diQFN+kFUwDlT3RyMGuxUJYz9LbEeIz3
n2KnAH9DAOTEEjp36faXSLx9slbuhLrcqmNrlednINdYaaSOjzGx2ro4dnBhMpEl9wKi5eRy0vpO
Xh+yknKiZDJvcW+RI7Q+bZGLiGDxPurvzRGH4R1gqzDwSjCTrj/ToF8PYtKPiIOjAFwkXsXU1kDH
GaRHNSxyrbhicb19CsSviUofMBN6mLniS74QWM06pRUJ2F6dVY9zCazDdmoPWhB2NrlmmUOsrqlV
eakS+viaMHzJxo7T/UmC20z9yeFAtliqBfvCWj0DNR0f8go7YyZOT1lPx0zN+uce+JauL9RDZjMV
MHflsVHCjSr350le8ZmlOR9L/GQNCsl1qw4+LhTf9MaFfc1QbzwregRwGW662OeHlNZSWWECtDCW
Ygd6kbBsyAHqxW7gTE6E34IqpvvI4tU/8z0fI37Pe5pbZVbhJ8wCf5QWDrLR+tSrdNZw2oIUBFu7
JTMn3qV8vg3u4UhTy4hDtmYpLYnwNNSF/47PQTg88bYi60YUnhGu5ZQ9TfeDw9w1JIGPPyeT+0D4
ge/sbqRZGv1wsjd6bvuyMpLvPOHnrDRvOCAi8MFXtFnWS0Vo4wxx1Tb9JYhM+xQx+Wj0KahGtW4U
ZX9Z/ainwDbi0shJtM/EP9kpknMskL02f9gXcujQIEEQePVkYW0ItqNyconIrFdE0+Hm8LBipY7j
y8MYDZI4sX+zbPLA8uR9QK87SL+Se8s2MtTDHlIHfOce91TIyA4RHfX1GWY3R/Jgg3RGYj/HjtsB
nRk+KH3uj+Do1dhbePVyAL3jzOVMhRRej4I33Uv3ENeVgOgNUpLhRDHr9Af2djG/XqdT1Xqs7yZf
TSoldGtYiGYUqUPcvjP+QEZ7hT95gCTF+dFmhl9ESlOETIvO46IsqiZC6OTKt2rXU7pQTyQmtIZx
O6bxQ1v+V4dXYhD99JhUZaFqt7ZJodZGfiqmqKh5PMOfLE/TLP9TLXrMihMHrHHlX8oDA6WxLiC7
5gncHt0Z45LBEte8E7gcEYozGvnlSTnioyPfyM6MCMSfGZozJfIugbkeEvamxsK/MYd1RG9a1z70
PcvqScOmIJ2lBG0Bc15ToUsxhLfhhXcHedMQn8NEQvS2Yr4n9L26hFH4M19genMSsRsSPDylDi/o
QBaw/Ue/IVNA9bKeiSel/yw2AEF79w6NHzN3MA8zax94PN2vc8/SwYHqxRXW4JwFqyIQEL+wVA0q
MIxzEaU+8sFeYJzzXfAeys32/7QW8MOi1v1ctWf4tXigWYqteqtEPa7vgqD2dcn9rRFR0swpHSSs
Oi+N4lBIqvF2E5VPHOUZ9CcD1YxK4MLnUF/Yp08a4QWSIPAc52omzTx39tjcgO5uN6dc8Bv/ZGdh
jFPmw3VZP4m+UdylWVl34tFdTodxt/HmgRT0IE8UvQKUvyzZFcvIpAl5eyMuuGfAyiZOh1NbLO4l
kkY4FVa+6y8l4lyIADH0Gq6xMLacocZg1eMD37vtaqVFFYyRp7wV3t185EJImveDSGJ1TB5dZ5ev
tWjzO8+SaJ1AVrKCADlFQJ6YiGO4ANlLTWhqGgIVxSHEspw0ca09k7ifFFDe3SSJPCyfPrA7QWzq
0ZI69BK+gMIJ2E7ybjojOW1MAs6CZReW49BiVR36wC09dbYEqKZS2CToWfihqaTyaqx8+fXcVBF8
63514lcNOE8Ryo48NnhCyU/NkvTYR/JDfEVJ6TvtfXrshmkfP0grNszoxceW87GYKE5+iY6dSzwf
yvoYuzjG2VND0eZGek9DrkSsmdHJb/3KNTrRzWaJHgPzomWb8I8aREuUBXpHut+cvMjVbsurvGfk
2wgmoUEVzr+qDVQrGQvagGGTew9mtzrc5AqaEQd4FVPB121LSMuOpS86DdYBVcZQLD/sj1TpX29C
GSwsPjUFqKfUa5o405V1B9g43re5vlxKq0ip9PSEFjs4mprDFhFgMqzz/mVspmUXNggTlp4nk8Vo
L1yILKb85HOGkta8MhocK57dof6fTe0ySjpg+QE+MKyshwSbBa2t53RWzctcAGeT2Bk+MbLq+lpC
b6EPJfv0duUa5ILdXM3sl288HqtOpef1X5jACMsegnUSaNNAxRH3EBMp8PzaoO7WQ43Rp7rb6lW7
14Fzs0M+xK/yK2slC76SzjJIXvL1nJFbKfEhngEHPPkFKTBiF5IlL1Acxkm39QocGR1MJm7qk1e3
/AZ7mZ81eUENvgPN9zQOMa1X3UBTfYT5cNt5KB9jtMPljq+3ZxjZNlD+TCR1n+I6sbeMtSiC3bS3
UYmeTb9O8mQixQDsG54nWS55LmhG5fS93qQCQzTDUWVvD4Uki57S97Ck5cqknIEvwMnnYTfledXy
npN7cklpRJCHl8Na75pB3paq9QjuZ4PU+44tvZZDkzYH9qgjReInLB9I+75nrd1zyaxJOg92Ztd0
tt8udp+hKwuz0MlegIHLU/5wcyBqZYJnollaC0f6Tv2ljKZomoe/R3pCJbmXdjCL8AUO7QYPp+Dl
ZeqCas0GTJ+RVJgvN3tHewzQ+7Ab+RSrXLev4+OWHSdkO9tEQ/+9sABj3v9qHl7JdNzhpsHF4jr9
oKrggxZu1Cxc8lA8Nwc42E4lmxD6m61K92laEfNE/gaw2mFyZyN0IjCqTiClRxxjSkT5WY9ePAtd
tZ9qywR3iZYm9iBtb3hPsg679lFP7xUTKkLbh6FIk0AJrubi6/1MG1Q2iFcA+bGPmw3/GSPNh+x3
/gN1lqAqK2U0/nJGrBAkVQt2OIlDs1HgYJbAHi5jO+eo1gqqi1+AK3VQ3rF4uJnkACUfa7rwFQmK
5IqJaAsS2DfNqWYsgFSH/97WhnjazCd4juOP1fVqE+tzgVuAjhayU7V75hpUfwdgdQ9XH/hR2qL5
QOl34ix4GGjcH1+gsdOSHubOIntbcgXaDT2iO8qUpgj6pyOheaTj41WBE2dcqsm8kJvnuzEIuSd0
q7DozdkQCmBKZlfuJF/6a0Ar3HWtBSv9asUhtrvST1oOrTNQ1P+68wlIizod1GbNl0xq1xaOvJxO
BLq3gg0NK7/XsOOg6g+DPMD/ukq+BoGo3y3rKZjTJeZ7f6gXU9cX/LMcnDDkVIEoe/O0ZvXp38xf
SekxbfiN0+QIa2TQJekE1ZNz6PYhQuCEd2rk8Rt+ICLh9kBKevmiD1jznXWP1lrl2b4/+uQzZecz
8v3rpQAuh5hZb2/UnhgR+WlANTz9W94YO3Qu1FBe6cGbO5vPc3ZKocippGGGningmbaGauqfkBL9
C3Aj9IGIi5OCRc/XzQcVwfZa9Elvch3/kkSv/Gjjss3jeJn+YND+6Se3pZhpkdmdiXTojWwrxKuJ
gJhEbgE/jy6Wzr2rTjp3gaHPkDJ61YfeaxiTvemfVetUJA33I+eJkRMMR5H5k5zVdF39itJnmb7Q
Jq+FyyueTXblOj3xkceZZzBs1xOwCYc8DntINcLHrdWnr0uACldNmARBftzXk3Bik3uwivGUt8Nq
uFe6fgAvMUBPoWdcQBhzl7hyHI7AEAPGJfUfrYi3OAmFh23g+cMJ/nWs2UMJ8Mpt1407WjE2sUhS
kTuvNNYDK++namqsAU8ioTIzDQWrp3XbrFtvp10QOBAZ9+HQk8lw4X9W0ubftsUg2eoyu+/0NodG
2CUtZCS16HKieLn25EDkE6RQ/gjRPs4ZT3OW/bYmiBci4uFIhgmusjZqI0sKClUBt3Am8+U47g87
9N6IM03dSx9P8OrhxZsOrhqrUEPXv+hJKiUT0MebwqUMLQFqLkiDUWzE4T6nPOJ2er//SrI86i77
/HyMG+Ind3e6o/Bu2/XoO2nUS5Ofjq6ZGW2NMu202SASaRR1ByO8tGxXOy83XXXhbyfzU/cZ8zTT
yBBhBsVc73jFLL3TJIleEku/C0b/c+QFgfN1GVD3GXPCwGtexjYuOOuDTzL649zLqDj3MRk8Dkh4
/1P3FhU0TD4vcb4CRhPRNgIntpeao5zSokSSJDkDnOGY3IWvy2cWfakJwKe/uU3fqwW8iHNQWg77
397IiFuS2bC8pu3HUAwx/yn4EIPZVIP6F+eEpC7k/C6cEuaahKYDfkI4U001r13b/wft999lvANa
7xAkHz+KK91B6H/cRWdDNQVJaK3aS7O6H45YXg59qRYDHRv89gL+X5xxM0lxFfdykScjKD6Qf1Sx
9IrxLx6x7dP6tsxdaE5xzdn+pt8dSoY1C3C2CdBM/roA3RwDvwPtKwpYyrZ4LYFa0hA0kH5wSNWb
E2Kpz7GgMYu0JNlLZIa91xAeP/LsHfzZFKNnnmW8JeMEPP/EgB9ydUzj0e4oMhfrX4/I9VkJclQ+
mD8AddhHDBEEs3NjWL61mgR1e4NzAoAgVKjMCIH77Ft4FDAje+9ZbWtTMzFIZGkQlGOXnab4nXFv
x/NGXAPGV/UoCFfyRy6MOdfQkJoO1K5cGtEadQ+BE3zaPl6mwC+Nw8tNh6jth1m/DLlC5Q9FrLhX
ZU7slvScvy0faF8fuywu+0QkUWyBUsOr+0kNZlzJhppMbh7xHiLY31s1xyM16CxO5IwioGb/2RyF
uXaD1GuxRelvniYxVgTOOwkbMyLRpDH7d+Nx0FtWfI2xNEAcSdocaSLq1s3HvV8mCrjaryK4p5fY
ZSXHlY5BUlYS+0dybSHeHC2XuU1TziK6oHjxs3yw7DXjUzkxeWM/Dy4tybGLzWvt+MPStOw57Wzf
C5I/EmZA9swOkdHqn7QN3ljeP6j1x11/d1MnOxKWEcCY4HVN830re7iq8QeTr53YttYzXJ7V60M3
RkXIMOxTUP+KCTP41hcnMLJS5ZRi4fdfYXCdVNGyP01E4WXL9d9glX/BQnFEAwXtTlWoxBS6FuCp
IUixQZSJyeiNZm0TLCPx9ykUCt5jgitlPoFi6yqzfCHbUcgXTOUrxQ+pVZ605js495ir7Vkqf+Q0
VdAd9HDz5sF6gpTNcEeamGS1ttHGyhc8lWtbgRzHdBJK6YKEQLOh6mA7Elxq7RmLKINeyLEUTAyD
81cNBRlA4rvDJLuC0EVHcEvaakoSFoIyP4pMlKu1wFHC30Qs7GSkPdE6tKEEPF7lWc9llKxhkpDx
cNDbVISvkZPNoqos/THe/bUrq0IIEjfw+LbpYO381iilqfMZbOQNH8H1zo7Ur2qr7/sSQ4gvuo1y
7JCPxx8FhMq7IUbugSswpgmOBCHIYKQVCZtKJGBSoxV7aJFcv5WMVE5fNr+xVya6DZRZCCf8oEHh
qC5XWeohdzyPz9YNabIiZDqyrFiELbUDHeSSzjU9625G/oRsmc4ewH3I0KwfxxEbGLwYSj1NDBdz
DUM2dWUamHYS7DJ8BDb2YKjMaidTpAgS+JAeEt9h0hTCoXO5wUkxLaJPXO7LbQSVPuwguob2+60n
c9itcUzhxO+CphvwNy8iF+fofRCqLD4N4M6Dxdb/p9zxnOCOZtlSpINF2HaAkPNAXEBBg/9IQFVh
nacCcd3fLQuMUEDELPz3dPwUSIsyJQSSmlJ0N44Qqa2lAAiGaHQm/Q2zh3VrkxpjMCA/xTB4L/fn
d5NBov6CwiiE/mQnLaHhz5JXQ7LPCZ9SKKcZ/SgTdW5cQ6y+L7Js3kqIaA7SyVcWXEl7OezfeLC5
SFCkxHY6x8GS8eNViLoPLsWq6ODFz/2Ums/mGbAPgsR68KlMQO9LtXC4qIBbmfaB3jCkni/OaZkQ
mSvLwId09ezYdwVm2xDwhPx49prSrhvTdjLNy6Km+8KV1e97+tT31uwSnL0EkFCBgQ9+Ku7FUKeu
088c65f3uYOawGOQC0tynlABLQpTesGojItpfBOBWfNXpi396lAeAyxRJcItdjwW1NBonMEY3AOh
SzDhoTJHJ3NJ6eosPgtQKzOyju8kA5WHzvXDkREaXe8G/Fwc7yt48fW1A9kBU131Rj+ZfEo4eXMc
5M9G2vHdgn4wqzn1jfMnMz0EBPR33z6cEd4qeNTq+K4LMr8INl/gjrZSyWzUTp8sZmPoFS3AO4Xp
lb73HxSo81sNfiBRHVPX92LhxXihHfE+iZALvS8bt4AXWhIRge962TwOm2QKE1dVGBsSQZ8AkPgQ
4rU097MhCKnC3rbbEnUnOEwn7tDi2EJ2GGTJa1WSOMiXqCA3Qevt1KIHAXSooX4w9nu07G0ZjyI7
8kgMR4s3+XfWyO+8RQWxG2WrjG78khfOEt85HXeuURqqaVpjZTNhr0rIdIxGgGFCb32JB9k1sIN4
IAnduY86OEaht1p4fxW/66mKgi6b7hMjri6VhZjUmTbxlmpXwW2Vxt/WEf7ttwwG14DD18eslAIK
AIeKbOqseYSyxMpFVIjlp4XXIBuoHJ4Io8b+TwyiwLVUE2Cs9IHVUxNDUHM6aUwnbraXs88xf+3I
RvjGXMwlpuHnV6vMC8lNQcnRfw6VssviE793lGgZCrlPChGwyZAHQTJTq7fFC8fj85bycONznwff
lQ8bARlF8XzMAOku1PsiOxOSJ9Ru2e1w9hhQuXSoYTwdPquVPHF1b4Y73rTUTNXKhGL6CRt5A8O/
RZ8LQyzn8FGH4yeNtv/He6a9SXRw/52BcNoQpxSkVU2Muov9RVDqBnu3OUA1Fmj4mJxDLx5tl9Oh
81Qa7LT8HF5g78jZ2rRhCOsWifg+GatEc+KUgyhK2O/bSZUCpfCLwQy7arY+Vq7VYlpXyOKY6Iye
BAIAq+HF1a6FJTLm0rc0DKrJpnU6/19ucT8VdeDEAKuIJ8htZRdZwAMt6DdmOnNxAKr4DNAngCV2
Ng7i/ht8qgF05mwjMEL2jbdXhBA+ghBW3tBsxRWikcRv7sw5JuJ8iWpvnPmp+aZ2AXmhvXp+beCA
WfNl3H//YOwTPqyH9FV93OPY5cCiAuzrwjD32SB8O12w1ZWtogTXxtrYouGG6OYuZmHkELv8mV2C
5xYk7wj+2HLeylIcH8/OeTjGjs2Pr/v/u63qeanUToxidgREptmFOrR9gI6t/5poUthLvDJwBfa3
JC8dwYhJ0oXDW+lhb/myhTfPrPOo4od/D6Eh28cqSEr/JpotEKSRAegNFjU+/ZVnnXF0jUQEj2Vc
3x+XYxSEacQNcLlqwnrW8pz3aPsHXZl8YaUaZUw+yYuB8iHRY3UPmnjP0J+3fIT8tRnOT0pxYR0E
BP8ZcmeF7XgHYavzS1w3IHG5kZ8wjFMS/T5orc7SBpa1n8z6WMxIGW4MrEbEFDjbKB2KXjTItQeK
QQAxXcEYFUNGMFH6k1LW/AotzNmcCC80FyirnY6htChHu8GXOCt3nEuPkXOy36aW/+UktCpbH26w
eY+BgoaeEP0oK+AHm2chGcwgvYswTiTxJ2zgSPwzEJQeT57MwsZhmG1E7b8H8TWyqBkZl6DqqU07
pmu0yDtLl5ti/hWVV/3NbWLrcHO690xm/sWYw5BOUT5o4csXZzpSWyDJLWWKWwxyp/s4w/yHPFwe
5nUk+rkLIVTy/8hTSLN1spOKCaKmgPJdu84MdHOyd9CecEfXyS5K20csmeTg9po/T8PGHzoa+Nm1
FN3dPapDr363N9K/MEKD0whZjZiTBoDZXsFldJmtzsxAoulonnFVgPWxvEXYl02yySxOvdjkAshs
d/4Q08jEd3mvyciLpKeFnuxdX+UTK8EOWAvKO4VsY1et2sJmDe2SIFBhJKebI8QA1g47P0FAYm6Y
DE0NP+QOW2vzAyn+hBHIkYEDc65nO6vvqYZ34auHY/PLMDN2M958SNYED215hkhmy6aD9TpdgSYT
6WCDqINaepbpA7O3hENftsmxn/8CqWS56WJuL2XiR3ubsISWPI5ojFBcv0cP/FYJEMpZZMD8B3oL
+ViR0Rz82w8i9ACYaDgqNByHrW0NJESu/55uZ12K6gT3FDfyDbOwrSYDTZeiih5+Sk4lZ2DLj06O
hs2SQSq0qxGj4Bx9mLS5Ti4Y2AQ8bgQSzSjWU7SzhBCz1TFwvunjYpKhuuAMCXM60redHWTPhM3c
VeI0LGR5eVF+cw+92BhO8/xLXwjpUqVvWIT7V+I7Znt/BN+ei+XgCYkR8ZPdM7GcxrVsFip0vDtP
r97VSHKdXE+/xSMy13HOMZ4G3nLOlSVYfDrCGjVTAsfxuQTZLkGQiJnpSygZukeIDTpt/4fQM0W1
z8lmWMZHB5NYu8vfvtWiI6XzfVxuhPWPPBhHTjYA6Q5EbiDHhF+hjDE6m7T8ZUARW4WMk+IybqkN
pIhX9R4vaGm17z6TgAhsqUKP45jLoTj+OVD4hicfeLyI01z3Cimu7+evPn7E5vy5BKAWyBRL7bcp
LIo7RufK5/M0U+QNCHmspRWtrKVHLSNQ+1xf7WsvD20P7a373EgR4b6IhvRFO0MN6RQzjT+bIiuw
p9zukL2keU5ekYLAvF8vcSsU6Ty60fKa5BGVHeNu8rwCUdXgpF/tt4EGj8+axDGOyMpr9PzfmzzB
M5JVKfGweZhag/mmy2GY44iLf713A66WcvnjBprc47IHaDN7I6EuG4moAbN9nd1VgeFmwcMldVRJ
ZrRf7FX04s1mpL8WIpdXPIEPH2L3YSYn7tJNDJvIWBlsKzWrZPTx8epK0rsUImNfwj8PW2Q8GSHL
iw2wLvoUhN3Nu3qkB7oV/VdxnbzS/jvJ3qqhhFJ46tl+aM6H0ej6d/9Uifd4UDejHSa4/sxmGTNc
HA3QX9IlzwhbPpHK9OpfrzyhwcqRQg3hlywzqWVnLCjlj9xHHrYYRCf9553ZMs5SMjTST5SXMnqU
tKEOvWeSq8UpcLgP7qz/kI0rFAaiKOBKxSYrwkF+sAOkiFuW13izJx3cRDmFx/ZlAL1Wv+J+rZPd
YBsQ2kFlO0NBhMeehg4MDXoO66Cs2rTHtpvsABzaV33HaaQZTQj7zn26wHaMTOQWEif/AsZhTfAl
GrtlEHeA+UIZPPKvZgCGZB1OOxulMefjoJO4sfVXhwWuly45Gw+IR7L8lWHUu6tagsSj/EiKH+zM
STUNkj3I5H5TAw5+ugFtwj5FOwBYBX4d2+jP3J4g0sktoNWBJum1ENDpZP2s+8bvYy0XMKmEUbVf
p54Y73AqvJPVJMUFHXZ6DGhxGzoNUsJ+ObISLnWZxLI6Jcxxidf21tauwtUXP9ABYecH/M82lCgZ
yOTbtxSn1Qv1WiFqJXrDiJ22VZLPkPteZaFJfu+zhtCXXXJbl45oIM4AbS+3+WWIdrFsIBPSPisJ
9AhWXTgsiw7o/9WkaSAb7umumNthl8bNeX9VZmRi8oSF6DwhrtTcf4JjEVG1YQttnZ2acm40r2jx
zQkgY1UiFh365dE5XdsKfhRTtAL/yoxdSU8kjAFWJyy3srf+LBJHcb6/EL1mSTSO8vBlW9x2YN1b
8XX7iY8k4h3N9amSE1/W6ws/DxkD6j5HvE4HHE/Zy47LhYnBJ667DXGAAhMVVQ8E3uSKD+8icLN+
6N0eB956lZV2w5uGt9irr0ehv/n3Ls7o4foyxbQHysktfAkO+wrwdIsNFAfqez5+rQLKVU+txRoC
005XVIX4Y2cFZPXTSowqGysUFX4sOpPKd01Gg6cmhwdmlvzyAvXS2R0XpHbfDwG0P2cECcGmPcWl
J1H5utIUppu1vkOxeo8pQF416mqb40OO8jQOYio9yA0s9AEsYu32+nN7dXNjt6iNF4P3n9QZRlRY
OZ7t5nNhHHHsfghOPp+Qkpw9nGijp8UgB428ndZz443R2Cuea9e8T1LwfSPMdHwCTS046LLdQg95
COp1a+js9Qdg04vr6yzvzAWvRqMf/cfBc8Jy2nTkF/wC3Y2g4JeQW9ajQCasijF9U8+Nbag/29jB
G3qDMTOsAnXrvDFMBNdDgj+vBVQwRT99wwfpsRQ4XEyrBbfEPZ6HkCH8KjWMMS0TSbR1lGBbUDGf
MJyN7C3aXIWdyGtY1w01GtW4TGptUdU9rNFFFdhJlCDLM5JtjJyXqc/2gZpmCcabhLc6EQQxkP30
quuzl9LTAyTxTOXy9OzTON0Jp3WoXwjNs+r2X2Q9Po15psI6dQvn0WkxvDJ1nzoF/oKGJdqmWusy
AAm8DPnEVEqTmau53giZZp47nFipdogmMCKcYZONL7RXTXtkweybCHalOCi2jPcriUjFB8n281kQ
U6gmk+C4wMjnYvKsZzao/asmMLmS16WsttlXGKDmFG70+8M28mDycWAjtK4pPZfiKUWDT/g5jLKk
tmMQnYOwKASIiaLbPrdkpws2Q/MdTxKqTPJ7UBjZQGvqBiJtU2gwmZbszoQCQ0vSYECizVtp6ZlK
kJeZMTDmxvI5FF2xsc64IYQZtoqbOQL5ev+2NYWQ5M+TPk48J7z6CR/t8A286IeWkVTp5CA3iKAa
Tg+6BTjS5JtsgcAcKy/gYQNzISnm7qpwbFJIFT8Pk78PTxQlIK8vOmtsscfmYIB0HuURBqoOQ9Ub
S9A++41F7qoCw1cW2Z2E5SFkaVOyhGGNVny3aeaA1rua8cmid08V++xVtsoVTsEyU2T4KhBij7al
3Kd3FLM+FVd3m0C/3HA6w5hhe0fPcSsFskFZT45BMoZPsqr1ToiJiEs7bPZh7wybgZSlGjK0zvQQ
WxuqZmJG8MGznWC22qb+Qd70br7S2wOwy7leCD5DfEhBdtx/2HJfv+1484U+zDnXe1+54zKFUB+A
1KGiT3zVzaY+W53drKWs0jcIp4vDyVu3qO3dKI9PC80fj6J5b7rml7PzEjRoSg+gIhc1Nd7F3fDx
Tu4SGSxCD1FElnf/66xKMSQVV9roBwqSjY8V0JqZexUy+Pe5wQPBiZR4DyHXT8ST+QPt/ohtyJYd
sf/fHaOUfADrm28UhXMX6t+dz8HfaER2Znq78SoesMlQucS8Jza7AXSO5IgLOuUhvYNIpmCG5EYU
XXu7RWMkhCuRPX0P7YNlFG9lsoWN6BUG3ciuEfPsqF588KawZAtCDBCjkC6IHzoW3X2nHWPKbN2y
j+OikpF5FYwEIDsAXpGC7+EW4L2eRElVsuWbW7gyzWgrRbCNpDUZifIGr8Q2xc9Fnd6n3v/YYiZs
ktk6/V6G3sfZCOvCYqI4PKf0I9K/sA9e3n/0/oPi4ydIUrKj6MKoHHrRe2YaVK+03cCLL/rIIX/5
/EPpg0YZJ4BW7kVKRvMXkSXmTrYN2/C15vTI5qzYRj/r57Idnh2HomOJXBu3wrsK4KKDybaI6RLe
VwRqxtBESbTjUnypap5bMb5FObLzWUl2EfOKv1dO5+mptokWgblwaOKfH2DIxVbiG4Lijal/vHU3
T2xZJmb23q2qgJL18yqDvPi3lfwP9ViiI0V3i/UhLp2JWzlFKhb8QUHmcoZ+BUivqWRJ3YLDUNIu
VEg88wLROwoNZdx8HOR3KiVFngzCAH92W32hxwO0gzhJQnYiRQa5gI34JPoD9MyqeTjkx3C+4ATt
3BW8/hG3ceSk4KbxbqVEKg2KWXbPTvBPVWx4gQXeUzcISGRETXdkHMZ24PDN1C+kOz+F7SjCtREq
Ni5Ufrh+O24ZyUbgzHFPfBBHehS4z4/01ySVSRpeiG5HztFdqLLmJWbpPgi2xmLauTrzUVT6p4l1
WEHPA0JwcZ8UdO9Z0c4IucBjPfbOOp9gB+msrmgWik4Veha7TIVtKmidYEDw2E4MniGS9y1g7eOF
z/fZ8azUEv9bl8G0F2Y73XD1oJoYcl3VcG37O2ES50cI//CZJv0RF+WhjniLunCDiqPduH7qBq+v
7v3PQEq8nIiBre4s7JmCVk22+aFv/80saoXjtem/itcmNlkPExOXmjBTIxVT7eSnxrGUQ61ipxzi
6YVEAeJuL96lerOv7QRSrfW9VNtxRcMYUE+kRDXZQXHJPM4OqINc2QlJjseZIMwUuzL3jKE4c31t
mzjUBHekW3aeKXBwYr8NNEaYaXVczfW8PNanv9qihoVvXEiQi45d1asy8Khku/9JwIxRxZD3giDE
xBizOZeoHb3/V4mkKx2X334z6of5IHrWyJru9UMEtiip5s08+P6/8Hl1s2EoCumM3exeNfbiKHos
NzYo7PSs4DdidnKS3ry8ud3ZOzwhUXMcwrZ+sH+6vrwATqC0oPzb6OKA1yaf+CV4JxEK+IKYUrCs
AaR6+Jyk+QZj/RBhCbZ68jPZKMiSa2w+llyiDEET6XVeDF+hRwtXpjeeoOtkUNOR1ipv3CE8KejR
O4t0sJWE+MdRI0muHnm5vOd45BqWOxUzSWDtP56k2vMudbBmEggK38MFWRbI7R/1o/kyM7ZLDXJc
qOSLhoE40lr4yoha20X22fy49cpD3WQmIQwxETtRxQwj09RVKWqj8Er8V7WssjRBCwObtJKWDYMC
NqlQ0YvVM5oCvwJDEvgNbd6PpxYk17M1mLd+4wvB1rVO0JE3vkFaSiMzqQsEeIxrHu/YkTlW9l6m
CKS23RrP9mh6zz1ZhvIIxMzH7X1u8mvDeOOXXcr9CMXtwv/RWd27g2lXI2dH7XjPZrDEIcLfjk+S
NieaztGuAKrVAJv2JTtMWt720JCyRkhtCgV23ap82Sdfkn+PnqxT4cHA7BoqDJnw9QFa0GsLB8Eq
dqIfQuhCVjAfMVREMPYy8u0KJu7GuHy+D3brjCTV5M3ld/H/GEjfOAFVr/7ELl8e4gJwHYG29GsC
lyWWwkKMB4+z7APdQe3bBEeczNaz7M8pPsTY+fdS9DfjlWafprsfPCkHVorcl1OLmP3VLAs5/T1E
REjoaDt5/12kVAAyVYR8AnmLAkzPrLDdvEHarbrJyKXIckNdp4cXulaeeweQQDmHNxIw+J0WZdKw
Bj7gJlzRDWnl0zGSGh7Cnm2OqEJgekleI2miiXP95K/o73tAuy8gm7YTlbfDLXBKGmu+/lggmBI5
scztgNYqPJzqcndq9KKSOwh+Qf+Q8rAi90X5AO0w2iTeSL0278+I1Rj5oYDPpsfdp+4hf7f9zTQA
5Hw+/giDLHDV3eHzj/RZfWTFg9SYV2B3ibBRnGGI6OOcqSUYghwDLFkuliWuBKsQFz1jVu298E31
rq48LmHuMS7bg4rHGlnrIBtOaWDlFvAUuKME81YNU1yUq3NG2wyjmqtQIl7I3r1ILEN/FQMQ9ST0
XEzv3YtSdyAqUOdOTnFtbEgQlUpK7Q+37atGbAw9gBvI/8P3D062N8dSamNDgsk3dLlGx6ltm2v4
Z3mz/U0uMvTd0UwbfUKD5i8X/9YurZDJtM/bqroAq/R6v/kMfMTCG8bJg+18s8rS90uYZYqwI0RB
ZLtHOIolnUOygJEqXd0lj2c3MOQ87eGxYbPQHatYpD68T+K9ECfrzNMa79L1LMhvT+pWhmuGE/VK
gF0+9dNhkMMbeIldLaWhiyOSZWKJo08oFgjOIcEHK9Y2qL8b3Nru4alhH4H5Zjh8pegvc6V2nDBq
yAMTiZs2qVKvVrmuy3lR71fCsOjZvV3tKWbedIqrtqj9UpXdvBLvB77kixXjq+7Lw5KybEJtIaKX
1Rbgqf4ykNTGwueX0GLoF5RLYW6GC8eeV5kFYpRhjEkVz2nnBgM3CjDCo923a614JzlaNGasl2Yo
3b7Szhcpr7PDOIsoJWosVySJjG6YFKgcVRNd1/WIsADXUPZYiwT+tBbFdpKD8MHwtkNYuSftKUOR
DaJNqgml7+Kp8njmVDb30Tswr8rHcq+zglNYetsKFAwnvKyzXHtGAlGY9BQiWsKNS2pQnscH8p96
6DMkl1BIR/oEW3rLEH0X2+IBATA5Dhd6v/fcfXvtLM4ABect+Jax1Qb3A+jmyoaAGYZuR8STu7QF
t455QFrUCPYxAEjCy0QMZvAfInuDzCGaJ1WLwz0RXsY5O49CkWUl35J/NLXBzw8GJxSD2qGtIxqH
sshZhOIIOfyUEYuMgF9qMEm5M69JrBXwgNi+UmVXMVjut6ix4lsfjpZO/iZa0+Z77LFyB7VCAams
AJUkAtqSlH4lnOdreiG8hUcLCbU4n+Ux/Ah0Skpgbl3p8gfMcI0pa2qBuuFb3Vg2243uuEFHRj42
QOg8gVzB5GgBQIAhErAn1TnEcNhuxC/fYDWdpEzf4+U1aLt2hpNsoaHwyoY/w7dnqnQqqds2hJxn
7P0yAuXrXWhk4GSb0gErw0f8HiB6qlVp/ShZ0mSYjW7RZEsffLeZPFGIrPnwxnUY2elBlN6UaDRX
pNCR7gMyo8c/OD1ZFiRlOSX5clBk7Gbb0IUCy2+dNLHRhF3CRWD7nmQwrg65x4epubWoZxGlTeQC
pm2G43OWyozjHcoduaLuM5d1QksoC5apaR1yl1lRon3mBGPKFyyAK3JJ4oZKnxoQSOESYaSJD+aV
/QqrCFaQbKCb9sksFZ93G3lq8HepwzqfZkdSRmjJO7NCnL+jLmN4ZbeNjLGDIzmj3SnLBwrM0qIr
OaIrkDsSIuHzve0WjckHVHc74gyQkyDxxHvePs3FSzg/Okvnf4kgxYqMcv5jxu7/OhXCCtLSlnQY
Uc+x23Xq07ctNYIsGV7BXACucqAbI0TGMEAyHSpMNwZZzcTKgQBFZmSGvIsRhGCCTdWru3cne77H
/4QLyS1kBNa8152dPZJbq0HvEueKyhveVj+bul85+/OIQ1gs6wLVOP1krnLLj7pp0vkDCXUjBbwK
LTm1wNudx0MtSGyW5bofwEftgS3DvzmeZPjSxULlCUJaKxfYZSdOJ8V0dYoPHLSq4ULOUtkbw9a4
h104GShZx5JgPhOer25RrZGnDSrd2tjrV8U8XbZjCQ+jJc4LmJ6i979bS4+SWXNsOUMJZMCPTpqL
lzC5+OF80OqbLvqzmiRfh8frbODbvl0Z4W+ocVfmeek0v+CnEJFP/DtTf8wPnb6JF57Aqg+xfJbH
8ndDGannqFw6KDc7Jry1otrDM/UKJKMftFJp1HUbzvncvpoXDOvemSLwePvM2736d4ydGL0bMu8F
vS0AwVReOnrEJoLlgCFZE5SGkkgZkim6iZ+rp1w4sWC/oGh2C8xsgRlAOa6+0i2wUhJw+xmpJHIC
SZ7ypWTjD8rEX3jOjyAHGw6CkA8CTgQ6F91QGpVAZQELAfO0AKzzOp9Wml+MjMY1LsQZmyqmd/ZA
fi4MBf8cAd90O/WrnokslUNsGost8Ss/+nu1tdxTMXurn8HNJbvbhey8HINXjp5ehtnqBr+pxwVH
VnfrF9kl3atB3vj1UECYgCL0MWELDfJYygNUJZ6h7JvEqdbnVGI4QsH9lWfcMvc6JnG54SHO2Dwc
cETeL4VUb6s5/lpmvwumfgSBp6IR1WKTKNm8IzvsCTZCVXMDEHwWK17KVB5rd8wIKUc8+chTwrfU
bNgmI6zWWwyg4P18EVSU3c3IJ+Sm56ZhPkeUvKLjxZPOgkvbij4yc/ya7OWxsv072pEzXYvh5EPR
1dvR/ShvsohidwlC0XfAVtkCk99Zbd1k+e39ZJihK1aezCeiF731U1qbhX1NEWFM5uUbBDc6vFrH
uR9P8oTUeq5KDTPcXjxqqM/Kyq7iP2OKZMUL4MmEv9pMu7gr+PlrPFbF6Ptx6wHyDeGSbbL64n03
/uC2jLuQvreQEy9NU3WPT0mff79LflbMVtqu8510DhqpGhhtLNOcLuMZDB2cRQ8YN8MWvztKo+86
Rv5nCz3D8OvseOlY6ZP8ws2XLwuyy2HiJn3mgjBfegv2iJhGF1cpSUZrR5D/+jyiQkmF+kaxNG06
Oepl2jOGAYL5spo6go3idQbsT8TDD8EOktGq9rXGD4Vm3PVHZezUhN2TvfYuzgdQE2bleChrlQYp
5lQ/70khzZEpS8rmnKLR8bDz6y42ylsy/+6ecO2Ztf2elP3JpqCOAvJ5DTBmSIuWLNfAjxgjkWKZ
cR2QQ7WMKwWMsqViwxmkwprd7T7F/vn4wvIsMM+rKxSCUBXIuYzCMaUPtEQWzYmAOdOgB//zKLEo
Rb/zntYSnCQlbNCGqHUwkBeWVC0AHXxLbNBC6mUSPFQ5I2wFNN2LC666m8qC60AkXZeUzb/bcn2Y
aN89MfFnqgMjGEkU9ZXHkAa6hHNdby4GGPQEIXpblp1wfVVe7IP26SVu4aZeBzvfShVQ0QNWkksT
GCCCMHwoSwKTQmmSGpGGzTtFoGcXthDVu64vc9lFvZdSfzFk3TRU91MOQcdiS88W4s0yG8kTfk/3
+f1OXCjAUmUD8egZ8n0/PHxZjSJ2UfNOJTWeZLAi3YIvYO9TxPqoqo3tYymNJTvmfaKjuq9pxIQw
fEeXjkTWuduPKeVGSVaCSoTRMUqZBUQZLwrMAtrZGUWUxNpIkV34bNxFz04JOJax9ZnapZfaU4rE
kcIQfv97C+i9vSHNTMSLILD1IK2zC+TI0/OlYs8LqJN44K8tTNML4JJjzr4yz8AWAz8ulAiMWOvM
fbPFSFkukFJXG2c1L+apVAM3vTrA80dgXCk2rJqoMNKO/r8j9pCrqwAMSPG0+VKclsaDzDIXE5mw
YjOTftFsf17/cFd+YTvdYLky5zIYgBOYFQAU4gGZHKbw42BWFBWSwIcKjxRvLTNW7tWHUk9qgV1v
T1cMJhcbuqHpcXwhvr14t8sFC1VK4QiEOytHCjpyNgUvV6B9m5+fxwAcsxXFxU4/hFC1O3UDwvDP
+GWD0ZbCMz7juqdcshFfqllTs9oyROFIahPafvAFEjHN1Zw30sZQT2HTEJPFOo2KlolNWEcFJFTg
LNZZ5pMvcynnSdwX8YxxkIIfn6TSyEueUaY6TpW9C/VoH9pwePpbir9/ktka3o8FQRdCmf0CEX3l
6RLpj3HjTephYAlVXeaV2dTmF8mCMcPVBBk+gqbKKe7layyIh6WjesHFWWRg6Hd1kgMErD/Y/Ett
GeZJOpn8KKEG1VcXVq4nHwGfhoQwEAtEHY7B9eWmvnzhVWwo9saN+j6HQkztTCVLEF62OX22wHAh
vd+TihhUQVlIDVLN2XA3o5NHwX7e1ITyn82xBaNffrHCti97Dtw21OylvglGCK5egzHJu6WriC17
6ODwG1QQRhw6DItQJ3t84R9Rs/Oat6wCSxarQiHKuvXMW8p8wd/1Zo0+qpyJaJ2a8SvMb6JecFi1
NbLivxOojUok0jSqU/rG7V2UfkTp4+1aR9KOHmYIGTebLvBQOEU/ucJPt3ATAH/WnIil4DOtbR4a
L5h3Ghl8AhMUnnlRPDyhjvpMECNaLofVig5jV1FMpRjxpzCAt8GwmPas3cZEA4pHFWr36jyutThV
O5tEOADUFKDuRKFFEtT5HOVeMEgPIuAd367BoHV4VUXzYgCPolbHSk3F0uHs3sSNS/oSUR75zi92
BGsFcwFZ8mLA9wgplG5m+JAH7BPn4AEFVkJXpt50yFIhlx1tPmYKGJ7iLXaVdywkqCBo+LbEOzEV
dzKAVoiA3VXq4GRUH4Qg2brWPmsBuy+QSNKvgbljfV9m2f3zmpmQjxGQCX26LEVMsIQBOMYKBl5Z
J75mozZeTlnG+CID8zyUbocTVBrbm/VcCcd5gY7/LFPbiTXlLDVMs05RWzu21Yz+dLuhf+bXYRcU
xsK4k/2Tyj9HpzfQdz8qzIJtvJ6FGQwALrqXyB7aNyzQXIk/bmNbzGCX7USBfeQ4aoUaASuteYFE
LhpvKd7iTJ4jBAaeBW+qoC61AWd4Uh/qW17A5PQLfryJokxbWahYbG7LqNW7pXt+NM9qzGAWBSFA
Z8+O+8bH6YKrcv7t1xg1FIU1wNIorKIJtgv8q0WzI0mNWfKjV7i/1v/8vPX+UA3h2Ti6Wxjim+pt
ARq43R1N0NrxX8F8RMnzzJfIq9Mst/y7PjtMDEjCmrLb3qXN+b/DK8Gkhhf0gv7Vb9TZCil3vc8A
XW/aztxdAZmVCtCRHdQhzMFlVUGgx43UdDFW9SArpzgJ+6G03/LKk3ITWgs69nLvlueB57M+6gyQ
YiPQ6wUAYU6poQ52V3rDNsRJK4b+nPeEtt3eJuoRQlExqQEV9ZqDs+c9zglLfq/nda2G3gsHYA5C
P7CZurMYRgZyLBFSVeR2pm0/lfqtA1hmoV5PapL87YnRB7UVs5KIseX17bfUMpNQ5xdJO9bLRBqq
qO5+1G1HlPV5XNUJhEhJfxH10YgTk3btKbhv96xtv3D0nNUBpIPvHCRmd8C1eIkJsWS2GGf48KVI
MDsqPaLAFpC6V9Jizl+OT7tPgzAZeonR+gFjKp/nviIvE7LYOHHx16TrWt5QDyb7B9pqPpUIr+nZ
fnC+akGsxj6CgOwSVMxZxKg+hE7UWzDnWzkiP5n3jFeitog8CDkcdOWJ9OXCyu8mRqZVpnZqdMtY
rxSC1ypmMlPtbcYaeFu8WlTz6HZQRC8Mhi7BKdDVn0pWS16LiTt/PCpcqzGWCxtEg+s5lqEJ5ob5
Mgwu+L1PUQZsRvXWKh6Sfs4F9H7/yVbyL3bt6IpKdCAMJuYTtfondFJOPZZM4ZugVsyObYJ7a0Fv
fw1TZXl0p17VTILeyXOqg00EM4hJ3WTvwCeeVZYUaLY8KDwSsSoM2r5CePEuqa9ygQFbrVe6PDWB
N6UKdfnOuPfB8CNFQ0CWL57BGaA+uRSUOjZbNL8/caskk/D3iii8oMqd8CYEqlgugvmxAinTiFHY
Sq+LorcyE3k0+gxL4yIt485pwwgKTz3NcKPgmzOPdh75L4bbJW9iy5EVnKbxxDOnsyve01pZPI9r
F/Frl5nCPHCmklmL53VNJGNa2d2iF0rRk1q/rtlqgGglVstjOmbuauH5B+wNpgRLmGA3Eqvxq9nc
YP/EbroOigA2qCGGqCbAn9/Oe3GjhNAgKGKDSaWs1UOX4vsxuCBQq0I6RTJgo7dYNE52G8n5aiOi
K2MtzcPXETpGOuNDG420ah3cXq4zJhdYpLCRM6bptejkAW9uYi1l/xl7jMxktwvuLHogclNQn8EZ
92U7Dcs6YImpOz9VJDtuV05wr90EvoQ0wFJlsk/zT7zCCDppWh1Tmsvvv8TbbNoXu54tirGYQU+A
epLGS6McHHMamglQvmcaQJrE2E/mzEOaxQgZbwg1mrn9coglJc+n4Wa9+CFlZrQKsK+a+EqPPhWT
M6/pEsR337mJe7W9Ewz37mBhDvna21EbdzMWZWBH97Q/sdtu84pgRF6OuRdCQ+lO6O+eIrziYXmz
qpYQEQgzncD7h7PdP+kNz12ogVeTwEzeytZ9EU0TeDkwxznQmY4vQFcSPiiNRj3X6OKfktb3h5qQ
75kB2JINrBgO3a+60U3KNkV0yDcY2zKf1D4mZ1WseqK2+J2EC6GwkJIDDizRH5gbE7u+k/wzwAh5
0kggV3H6TH8AIGawpTzlSwaXSz6QTXdRKqgr0Kt4tj8UZlbsDaxLYjsZVi5YMuT0WIP9O8d7/Rhr
Pc6oSzP3EbOu3JgvIOQnNQE2OC6WDINtokpQ0uFXpoLLKWg2ijQBWiy9EUWz7bx7OfS7Zk3+UUX/
ymr6K93xDrdYom9VIC/rYX+eBXch29Kgi2O+81DP7ML7PPwU/p7kTlP26GRrYbKEQU3z9SLaSzjg
tNoP+l0uwsa2+0T9UcMQ3ODPrBLWZuDr0vdjdAcNwd0slMVcLjz5sctkB8yxmoUrCU0PBHZABiS6
HavnHzyOkkNrD4qQp4bYYQcxXL6HGRQLe+YF+SVqBuw7kdTWTnsMUHYGmQtgpnitwJJ4sngb6KoU
edJzuQ4b9E4BGDKphL0h6lBs1m58AE+LZi+XNvHk1AZlhA0KQuhQxB4qz4A79yVz/Cc4bxa5gJ5D
woYEshf1/aRCiSYs1TcWoZfwH5xJ05RzxBhLb3PuAgX99bTouehmRvpu3MVtOwKZB34qBbcUK6l2
Wd6M6cWgULwjEWDR3+gv4Pj/zpE5asG+GNTij2d+AM1xBiJK7/eY1Qzm3OBOPmxPY9MtNl8NQDmD
LKor6l4VQ346L1WWtEekj6yOt/uyAsFzRj53LFv3bGr4ebpPn7GLx8Gllf55XJD0NPR5ik6zhhdx
HXj9TvzcR8ua68wO7G6VupBujEEfUvbKKII/D2EZzRTAgZdq/IaeTedgNShJIjlQg8FchciHTIl9
DJolzU2MmJg5BNRSFAjF5VqVGS+4OARvfQQkW9U3OWQN+9A154J3GLN1exWkUFBDDynbO8id0oe6
U/agFeBohETwz2E4G1g7ezlerpRy3J6Slk7CI94FcEzAGxlXgaPBnZl7dD6Ubzo1Oj343UKCEsh8
vS42SWHkU+tbS88BJ+r8rAPMijfgX3LgP+pJgicoDrUjg8dESwHXDEcMoQ4/9Q/c+bayZ/etfRq/
UVQLMvN1VgaI8RpiBTuOlRAnhhBfye2kZf0G2L6EOvZXibgy2Kk5NQ0JtL95vR0vBU5PhEb5h/l9
K7/UrjvY0xCeRlDu5Cn7KTUKX67rygxRWEVFQ0X1sb1F49jOdqphLVH5CsoB4mqF4qN4UZoi+h6e
+lwVLMDurWAWTcZtcnUYzAQZpNEkOfHhLY0tUbNy52AYFbo7Rzi9adoe4b+DLnSRjbBMDGV0xNES
3Sm3RUSNoIQQOZlhEdmD0ZyoRORIKRO75661pjD/LBb8EiasaYM4tBnVSUnWkEBaYWyZiE8+PZBB
1GxghMnbksWyA3p467fmUdYxphvLfRO9ItbGQjClqYIXgrYMFvruCdT6BBKowsCzwpxcZ7pASu0B
CyCdBcZ8gLrV5Yg9mpQQagZZCY7E0x4xyhQt8upSotdIjCAnHSnZm35E2ZqKlKFX/xr0s3nHGNoC
nnL+3PU6++BZcHKLAzf6EBsoBSxVgbXyxR8ghwxAKNMGRFcPqVFiNVAAM8UMjB7XPRDLzYitW+NH
z6DhTmMo9lNNT9V+E90in2f7cd+sqDq8dRsn9sYQf0AcIP8LhSLD2kDpPfjkpvrXG6hr49l3q29s
V6M207pvRctKRaK1iDWf2NnYZKiKYiuVmy+M1cl46mYHsHp8cqYil2Mnkv5UajcyZ0/iweug7/kn
f8f6sCid2QhYwkwRcNhDaIzs7Xyc0tv1pyL/drZgSONHzTnKPGi424pLGgxjbUgZjoBZcZMHOffg
HQfL+W30OBfjq82t0pH0nESHvJVbxRZmnSh0+N285rVuJ9VHrjiafBqwxDmOJGQLFWTbLpElq2kk
KOQdTPCxXL9cj3WXUTRfsu17l+0wPICDYhn7odK2iE1rH7etjbIyEGh1i9Mkj5ZfUx96xsfs+hNw
WsZ6y188x6i08z7XXAFqbxKLTd/2f8HxuiIGccf9+ZYaLpN8S2tMln+fP8mariq/vMua4dqIiREW
cPHIqdLJBIcuLPCnUI2kftwSF98ZRLoSF3OpNDOf1hoMw11pnCDIGeyv/4iIaxK0f5gkLegdaorK
0BZl1p6y2HjHIyiCnuwavWbcewz0A6wBFm++Fl2KHb5bPHAPfemLJ+d6ToW4UE88qXmVSUgZTyKP
QABwPLt7VWWV1Y/BlIg46FijTMNEeyPmT6FgJN3LyXKOSc07KrwUCFdtY09DFeQZCg+2H2TYJLvr
i3VUntBxD+IkEpnThVWhIi5QFtAORxF6QMrJ7sx8NjEYOSp78YYhlRik3lHf0zQQfkI70xoqQSN0
zT/kyay/7ZogciA9MQtPO3GwON4EtmTSUWVwDiAll97D1tVwCAmy4yclnKt+XKzuELbO+ciTOse0
662cTjl9L9pqH91tsH6nLXdT2Alpht0PrdH7vB+s4/1HS0MVUoKhRb0PCPVJb6eu2MRExJQYxVWV
KhLfqsY2x/AHigOtLRtUAWhxG1ZXF8tYfJONREURrnICp1k0DkowHxL23+q01GF/7z8HL1ZPVatk
TJn6EI6As1cMufqBseI5bIeVrZvqictBTrj0Pf/0a42DdQc6ou1k6ZewJC7Hk5khoAyGbOYBzUhJ
JRSQoqOM9wJAiowNkmwsujiEd3phtgxKVBIYMOCLylhwjBYP8xGiW09OKEWzrj5EH5yBv80KO8Aq
92FpUm63lNHJ+vA2w9WxlwdQ8we33NOpnT/P/N6cTLujHJw+4TjHaIFWbX5u0yhZjvCuNWQHz4t5
z3heji8ucI6j2Mw2fcMQkRykUGlT9pQiQUavtmzz18ggGMbMEs3ofa5Niq+eGgN0iBz/OJxBTsUa
2gmwSLfXD3eLG9wIJXjSZ15hPKNfGe1b1a1K4cb4IIPjkQ+wylljxfAsWPnrAD6guIsUViuWZaus
zaz44U1GnozYCcMmQoOF6YaNT5CDTSAjhuPmxqvehbp067FXlS7y/eKll95rc5qaBN5qM5l54TcR
5f/amf9p60KZwwB51e3kg0I55O5tqSctjarZg2z51wqX3J3Q7cZPjU+VhZK829oTEMy4u7UMghj5
Wvp9BcGLFDPif3fGkJvU0VVoc1+Bq5fVpRnM/hCgzgxGiJJCTiGkzX2SzqenAuQAFk+gpif79Buz
HY3JGPWihVRpqp2Xd0/Zre2WCvHK2q2BGVNfLfdk8AiiO0p6NkRf1u6+HK1ao4AizBKTHVNXGaQk
gtug3C3vewoF0REI4lbwuvV+hWQGj0aBA77Lz9CcybcAoimjvC5akERF4pO2aMpQee5odFewCnb9
VPROOVF7vXAjgnxOAzl7ssQmaNzk4P5wLLJkuC8zTFhFX8VcTmepD8iUpsCdddL+eY6A2ZfUqbVv
LX/PncLfd5FVHLwnY64DkWpNbb3XlQ1v4pJtNhdcctmrQuRQ+UOFkk03OV3JjkhFslTL5WcX9cH4
fhqv46lQnFBOPH8XoQP5alqZ9fBp8V6J/3B1bTOXSXDsQ6NT2lZEqAZcBQVLZwZXcNHXO9Lzbjxr
1x0fXa8cPIBIEWM4tUFWl0ycxOKsvlQhybt8b0eW6bkrOA5W/gKn8abpfsNhfNVHMV5Wj8xmqmL2
43C/E5YnmIg4U/kZCsE4GPQduvARoXZA9Izp/K7yZ3uJfTtr04GOd3Gdy/v1NUKOZuDMdcwrsflT
IxGEN+o4wriN4/RQPio9wtAqfTK/n+xq0i8kC843ALJUzQu3CE6E1Mj3lxqtKXegfpzr+tb9tWKG
1QKH8S0yUgHuE/c+Q5MfYiTKhjF1Z6CFypamIipMRutuhw5vwElc2ZD1xyczeDeuLjxwFsUtyzV2
5iSWFqavjHieh4NuwcZ1Hxq0bQXvDFqEIL9IGaG26HjAU/IUpUuTnXJbuKQ3I0UaQjyjFESmmlZ/
hE+FA5kUvi+ENQ5hU8mToBEbE1ewgh365itxZRtQvvL7f2OoSQxYBpRXo6Dr1Zfk0T/15gJ+vhJ2
OQGxFjDK3DTdWDyAiggrS6/XlQ9/iUFvW4DebVAOkJyBpwBAjBRRRq2LOlW+3HHsrj+Sz0i6N+Pp
LzkDsO9p0WyWaR51yVYzs5Hcuzp/z7ywOumYhBPDsYxOWqWml0UtmM7mKn+1ctZKAzT2GwMc114A
QHqVcHuwglfhCuPHX2kc+Egr4h5aF/ImoW6oKGrntCoCrk5az8G1dxV4XyYOQxgczM+r6L333hMv
ZfEH74kKhQ4w/J5bRiJJu/9n70OkbD0G81uRpisBaimoyOK3SzBGhPXj9WJX4S0zHrmouxzgC99x
ToQTxnRZ43nrTbiM+IMjX0RD/fBax7DGKdJT+ot/69ohJA0Kc7WkSl4FX27+53YE4KjDk8350QO0
oVCl7Bd2tvcd6UeRw5Jk17iPAytMgk7TVcvkhmCY0ZPdDoTcQy9rHxX5UT7efxObZrePsH77mtgP
CmJrmNwuUKaq4QICYb35FwVNC/XoyOmBT7hkrnl1IADmogP9eSamiQhvzwCJUTJhbVfBNP8BlJHB
LYRk3Q2pThra4tyN33kEw9usPvAzqyr+h4Upfif+Hp5y4NdtQLBFbpM6v0i+1clJ8xthY+Op4JGY
yIo9j+inMwE0thX6FNB1MJzrcJlsuHTiAwcx1wbVTIp3K9B7HDR+/shZLFLMpsmq0z+hnOwlygOQ
sVnuO/rA95Ddu21imyhnKGG0Yl5Ty3yTi35LItx/15ugzxI9MKRFS+ePxAZUpYuH/K3UnGj1cYK0
0jxdaIi3pzRAHpi60h+oP3ZohLnVk/9r2CBFPB0th9QQXkcVoFdpCDUV9qFvrRz8wBdWE5DaUROD
xUa0e0arOa5sC5saX3ZhZqslMt75MHB+WrMiPhmMNIRfqYevHqI35hWJWq4G2KyH/mCYPXx8aeNL
e2jpEKGovFXzVVRtegz2DXPxiI/hCYoMR+rMpSjSQ6RRycOwzJP01dPoI5CYGZQhQk7k8LSqSX5i
18mvNx/5x+s8AGWPs7fn3sCnDSYzGIyP5BDH/Iq3l59If+us11nZ0CNJFeASr739k5vshTFBkSDF
NZJHr6R61XUUqM//6SQh4rX/L2f+4mY/duMJM5l723U2ZTHSUP8TtUiG8wySU1DMkGPxZpvc7ad+
5wQMeu3vvxz1io1VXIXyNq7lk3FhOtjYZgGd+6BXFph4VtD5atGdr/aitd6Epq0T+iMUz+G0KMCt
OrQSF2Tii0juWVP5c+jdAG3k1UmXxIS/0X/IZc+H1wUI0b99YzsmCMMzFuaTicsvxJSS84C8coLc
iP7Ocv2y1u2um/060ZyoolAVn+R2mCEgcV5rvCYE1ThODCYl1iZ/u7A0VAmyoj+DRG9FmscYSwbv
VXoxGoGBTpk5+ni7GzwAWc0Ch3+0o2Uim9Luecr62sbl4cV3tqBVt7srx7r/duHhOFkWlEZt1tk3
MQm/QAQks9TrCPo+Htiie8rAdKUc/H20NjM6HCcM0+Oku2p0vwcUrKSGjBY4E8mlLcJ1l+dq9bFX
K8LArIaZEgfD/RexJ7OmC8QAfTbogpW4YX1DQ3pTACjMz3P/358gkmORZnlE1B7Ff+lNVrTFcjGo
duqK4vDuhVOF5J9FqHbObj3W7BgvGYIOuV4yJEKdUwA4lfkTpxQSRJFoCRUqsC9YSkaPjt8WYFID
quj6iVu2p8wmuCU3oRgzV7DbdfjOFkKBEGLwCVj/ciZy7sPN/Q2+bS5RB0D5hGIyMcime/wiyWLB
BgUCer/LalgeYBxkdy1awv4GfQFIPE4kq+pXcbp51eVwHlA089XGCHtwdD7q+AKF3ggVL7IPMCDT
wdGotppYYwvCi9U6Otu1TdKCztB252k0XezJE0zZP6Y9lIoOvoyODQQM+lX7oM9+8iQTADYw4xB0
ILnJozFnMbSPJWY592K3A+8CaLaJCX4XoT5Ex08JSw7qRRoVwTHvsyh0y4ssOK2GwWiHun/ivFiG
wsfMcE0gy85D6Zi53qIXITFOnu2aQhanaxlM7YEbDQjcf/FHA4mDHK09f05cZoxWng6QXD50ZyNx
7V4JGR93Vl47JUfteuvNLqC7HHmvXcyAl63zk5pq4GlAZ3Gsb72/E92gL/AiqhXQRKLcz07PqxV2
USb3yJOb5rikmkQODQXfM366ics8FI8UWQg7IQJNhxKHCSVNr2y8ZHnDPPBMkPfdPCGK3vN5uIzs
ClDAkxOLLlWeae2+dBWiAApZn1Z+DVK9PcBCoRimmUxpFKoXUZ1AQQEdY0k4tNE0mnc6Vig3deZg
TcjwtJR354cF34rwqbwJ97Y/kRCMkzfK/e07DxOJlL3lStQgbg2FZpXi5Q9G2o1FY4RNF4LipBil
RBPmOS/qwZ1dwqYxsNG6Zkfxhgtrz73eqBywThbApMloH2ups9a9ByuwytXyDfOfYUALXKOweaep
VJa9cCJJtiHUxxXBjDw0CFQ58E5BS8MvVE4grdzdahKkWXkZ4ys1ewFZCZqU0WxkGX8tuRV/Zno+
+rhEdLlY2y+V9zZ9kQoAasLx0strPa5ogtp/MecgQneANC8HDZOdua9WjtVEyDSNqSGFNGMXUsvL
vOa4PugDyd1sGP9dLX6OEuDm8dRqlNvGxA0pPcW8av6+di3+WaBhcFPoNozckY/n96fYV7z3hyX9
jW44P3RPqrzIKSYrB5hkfI+aUrEdeOCeMQAJ6gzJ3k+wMS4K0WOu8IHGAwgQY5d7f0nMmsJW0A2E
Ulm0HJON3AXCpesIAMxnXf17QUVjHm7cvWgWoxEPJA5o0AH5/OeIsLP4jbRDx7xyjGnueF0ML3B+
cy7WIe//olr/xntHgsAFdgtvQq8Oex7s2YtMgENvQgxUenWia7SDgz7gUCkFIndBQXuGSvudreUg
+D559/l743vMeJUEyhmZQYqB0xuVb4YtRcIS31U3082+SAtLU35/l8/k/zJxHdZuIs+ADNVIXVqf
qTv1H+/PKZkOpgFfpwuiLlPmsx3ZHXeB0d4r/3NmGXxkjG3WKb6xIIWQrhAXurgtuNIbxIYipUls
2V/InqOIpn6v8GCpzh091unMgIJqyg24Y36qYLcY9lLDt4YkSVUZMLIlbAvyh1wrb7EtpvIGrbB+
zaAvOtxxciL4ErsxgMGbyDVk090Y0BbLZOMM8LOJqY0Fv+MimjQTLA4kzworUaeC0SSHN5Ezv5py
nHNstJnxjsosTp2SQKrLjE1AbLo7nP6TS2FhKwPZCjyQ0G12ey8zpTRfJXY8W2AhWZFWu7fJoHbg
pi9Ug6Oa1pbFG1Ubl8YiZGKEdpKjW6/GTLnNTY9+H4nbtvq5fpz2EKgR+oaY85MmX7FH49hVlL7p
6YTHOT0foxj7yQpTmGXosP/Y4WLSDo1/rP6ZnOrGx1bHBle6zmP2BMCHqcR0720vnULBWBKDxH71
sQ2jFnjnzBM9vtDX1Xc88h1GZWHjMo3ASrVf6ACH0nez/38hKFvz9zMnr+QRQ+2tTR23Kc8RZcsS
7MM61/wFniie3/Ge4R1GklLUUOAGmBctAns7lh1m8/43EJnHvcmSwadr4EMDbZQbc4qhdRhyvq8y
tf5PzglPWeTXLSbQWemSyEeaWo4TNs+VHx0+9qzURSMbBSsj5naar6UzQh5HuronovHTNNLbfQEC
N9k7Mx4sJIH5XCuxOimNGS93yA1NADum3VgQC9hrrLGTC9SfofndVwTPcPu04hWMnVcwM82XuYDf
fdpxT90FRO9x+Cxxdh/NC66NbQWkT8hUFMYZMyEtjEtHQqKcJ3UVjh9DDemW00iRkmx1/qQplONI
kdL+CQ37QnZivj9ALjWJMaAEcvaJSNX813gktqQ7neaAmqpUK8vSYt+pkdS0k3nfrlUAevTAKgct
jXbQjw3BVAWNKanpk1ixZSRDW7DyhcLAqs+bFJAUnj6brRgSYa7A9HGy6X0awov3gz7ij2fPDPzV
UTyrZ4yz5daXeDS80t4gAb145CYLukyvVAX9AeoZWYOEBf6AdOIkTJZdIg9lQELPIbQW4RvOjL2x
0FLqdEfcWv+2GgNv7pHsGf/+I0UQ4Z/3dwrjgvJeMHZeqmNt8UtG9J5biBO/NSJdjLQj47SuZ1SK
ILqaa6h5Foby2WWFUQU7n0LJiP8G2nrcevzZo2dHNqG2UhHhf0bzjBGkqN6hPoFfZSzPYiJHEGrK
6NqWXRhcAC9l/+bILY2XMYX1yo31FvC2slIypuXqjpoCc8cyZ3rdJ7m57H2tbSntCgOhb02ZMPdL
/rdLzzIpBNQqcxNjAjteC2bcEIuDVwnQcRAc8GWl/bCP1sXoiI807Pugd1JwKth2XVHp4shHp7zJ
4mlpc6hXEbCtRGmrtizYhLmFzXLQXv/zP0oUwozvfh7iwHRxbf/3EvmPuoksZW9suubzWMUHROvX
zkmMll2bVo3tRI0qfjkG8s9WdurLfofW7oPPW6v2wel9FpP9EJRsugVVK4zENOYoOCi2BQbjsyZz
GNVj3XhzUJaCaj2YJsJfvD1NFj/3q1MEAWCcRN+3hUBoYvdO+pETZqhisTfcEmNqkjb6M/SgOLVB
pZ6inzrePJQRwDsJopJckezuZrGIr6auK5GVEcOLVBCuB79MTwNdUECpGRFcbLNg3v2QY+tg9S/9
7aTRpevDTaMOfr2KPiRaAfbr6lVUhjEs8idcCiwS9a++zF6mOucTRvFv3uA5uFIwwksalZsEJuJ1
ninmh4byckoyGJwkzIQttEHIJUrLAj7QbCrPYfPwP1V6Ha7KGQ7bnEQ1QLHWRK3nsuiVnOYMMQwp
EqRcIFxZYRWehJ8v1V854rxd8q5NkioUhV93HVTq8ha4HVOlRGaq+SfKz+iDONyX67Avip9J+jl+
Iek1v88h/yE92QJQ1TtaDLbiD05iW0CkYrOfjfHxVqBsBXfye1mLdPcwCdGp0ftZtFkr8tUOYSYB
YsmhIU3yWc49OxRhrdlGbIV6sMLrsS0PYQZfspZx7bkd333jlLTxBNqJlHy0ckMhQFut7HtPdMtG
a82z9g2t+0QjLODEZ2zEa9wfnWYrGeyoDNt7l3GaGySWAtUsS03IZriMgfuALrderTBsFI7gQjjd
wz3Ob0n/ox/NYHmJB51DDKB0rNLjPfAWYFsgEHhbqV9iEKbUAPFUncq5mwfAQQGeT/LRQ/JNEpcn
HyU9erNJ09QH6jn86aXgxbIvucm/QKjKhoo06WbCrDBtiptUhTfN+HY6y8VykbsQFTZ6o5w5bwrI
pmVlLKlR+0n2D3GkBv5OfNIPIrPGAHOmrR7PHPtEGEqaDHFE8fpbgLh59KQNr8anGC2LyBAiA43o
DoDaUoqLpi8vnQGNUaB9sy8Xn6mpDg4gqLSU3M7LRNMXXW+dPhgpeJqTVDSc4vNltRKHVjsfBJ82
uKdzgpBa97x4JrR3LPE+9Jb2W10fpae+zYrKNOzJGpbrrZmTwxas2iPz8q7aw52XRMRAzbsGnBiA
TPoAKYgkznT07QnfH+XROycT+t76cnVEyWfZrBDvMVWPqrjtHKIyjLR4CGqmCEflCQ7MMynoGB8n
EW0Mi00es4iErj+56SfA2hMGpg6LUN+vqGULICSVsUWwTYoNMxR+TkibT7iwifpL6VzYPLXVuP18
dzZXAWxTKpsfZL964m/aPxPrPeOloMF9qve3CgYcEZZnEXdJz69PjfagpISPstdN8xhi5wY5ROWU
+QwT+s+yiJ5RzwTV5PmKIHpYgYkQyLCjXC9gAYjARGxSiWkljEAar06+3dibTDvm8MRFtTHEXKI9
PxMxIGY7kNk5qtzVEEX4U/EPReQJuTr1ruaSzo8BthY4K6iF6OisBCPhFWKQbQW2qMSO6DagxiAs
qx19TbuR37gWTmwHO1NpSWcu0h+HP3Ad1RggKEEqut9tiroW8jEg6y2bLo4su8kknGkuVNgtLE+8
r1Jbs3AcQfqeon8GAG4DAH8AmIgt7FKRZ4v7AVPovgu7xoHEfRhhOnVheR/IR8YZOBWfB5Wcqz3i
3dGmiENRqy+qL1Mm5KW7Xr9REAXP/wSJSXXTQJfXktCax1Cjv8p6FssDrdXtMnXYBZoxiGTuxj0K
xrKIunH3emSmrALUfN/uG65l6bvV0CWaNaw6e/zkc12I9pBV6Ci/N0OLDl+XDC9x7VrQ1sYapSq3
/omWCa00oAbMhNgQkWfRdxJLvry5V0y5obrKPjBy6Gd9u+xLdKNaGow38ufdg1uYMxzl+dpkKb66
gszfdrQwjvh8GQUEJRoy3rmkcn/pEbVZYKhd12ofllQzTpqRO2mzMecFmPgZC9NvvqUOwAnmSgrq
ZB4drTxXO91aZ4l6yX7R00lMy8I8I5Ea7A4PIU0dCuxuuxVn3iJSwfMZ8dXbYRpcr0HojXBpkR9A
JqHL/XrmS/Gk2DJ5ZV9BOUd91dMq9jEoTsNfdheNDWgGNHDOs4aS0m6sY/gaD1lKRfISXclO4m7U
KHIdS48ToWKb0I9dRLeI7TBvPPgegB4C1XF0Bn7ytJywQTYjpEfS8ARkBqZmODkXbkOL9lzOu+i7
oe3f9c8JX8ai9crhIKrontJJq3T0Y7qq4TKSyqZA/Fstc6AWdvZwV2Z5QVPvVbvwGTf9kbapBpRT
Z1lTrFZtNGS0FyJldq3yAI2MKcv5c3+HQAT5XS4kp5quVsroJZSIc3EPDGbGFXfbYd8kqKP7EKut
OE+bSGaYSrg9gPo19VUTLqEkNvNmBLV9B7K5uvWb5KS7mv72QgLVh2+xnMb1S5b+80id94mEdPUF
I6pc9GGsiwRkiU5Njq+CXv0m6F4G5xEwbbl2DjtKCsKcgBT12elPirjL6xbzpgI80QlJk4iGGqHc
0PFVgd6NtY6LvyjjFBkajHDgQgqiGrZBzwHA/qMKxrEcJywd06U+TOJXVHgHIClnYq44xIuhKJB/
A4a9V6/njbMmE45dLmv0ii55gewH0+aXD9KZaRKpJGi7Aw9TyEKRLjA1xA1II9DxJ4zyMds2gZvx
sw9+IFfgROnk8YtmU4qdQ7DBRhGnygtBg/m/nXpWowvCMs786OXt07g3szYMYgzLnuM5NodXg1NK
YvEwX8zFacK+FeCTF5fiCdn4GpIJL1NBQNNe27ecME0g/MBKsHynMiE6dPmsYMrWZhNDj/jWRemg
7y/d3fDSJ+IjUw3cUz9L2nifbgxjxTzRKz2ijhnTKkKSbXk5EBrtK6x3x9iWBz714AYCgRzL7N8C
AHFTv44iuMbVq6qYsNNEE1eaTdOs2bawOwBcOvzIhiYbasckk1/M8XMFSgGZTdVyVf+wZxVXbk0P
8j+1/kkbkWjZOvjPHERQYMm+jnJPXhdr8Jg09jh/QqEqMXry8msjsy0E3X7oPS4v1SdBrLiStAzE
5OT0hsD1rUa6WFBjL4yKLwkS4EwIVnsV57svp3yPcJQstTqfZGxG2BI8agPrQVtXxSDETIRwgEHN
jnhSPo6SuUiadx2yQJaFHlm76NmZ6ycnhG5JYT1AOcuLeF5KKR+Uj+Lvruxq5ayYuUE88za9NnAN
rqyJAOX/X8k8a+g4iDVFfNcobwrj/FdpWs/DBofrdPcV1RG2KNf9ucoPABicEq9uYOTllOhJ01h9
c5FQEv5sRAhtFgXakI73/QFgiCwmbncbdlwQiqOyGK5h0FfqQggJrCujmjJky5CfADG9G4Y952tt
4kq2x3SDtP55tX/FmfIA9Nt/zhB0QcCql3efymbFCaiIhOpms1nWVJSUfYK0cxngWSWYz3jMl5os
R0bN1ahUsBYieAaanGmpcF2fF4Fr/DbW9u9CbBrtCZwxLh3OleAaGKpWVRMFjoq2e5930tyWEJ17
w8XvdPQRwZUfOcpff4Yv2jM4Pm7YMQNMojoMHUjRRBUVcIgpqmfrzquexHM9u948QLjXrJCBJxiV
YoaAVzka4B2S0rZMaRqdSoimRn3gzlKn6DPixJWhuR4JxIfksgzEngW3aIiTC7TOQAUTAIEHBou4
V1wGSdeSsWZMrCgrUTqoCl+TTpvWbjPi0RtQVUaQ/dLLLr81afKInPLueT8sxlHdxTlB61CcwFID
TdXFOwNrXZJ8/PNjbF3+DeRSL9R7FtB253P7/NpKV+ZW9NlSHwF+hYwpdqHKsptDFQSrE5vQnGFg
7xdREauWtHOrBhDUZ4j4m82jZI6ejhxDGJZqtv2Dx70a7UArqIEAz1gN3y9VMKyvX2hPPitUltoa
MEYjYYW/oHWCXFHYNnTPaAokRcLYTiZauVapCNpmsWPPbcPU/ejr7Fe+CvjrhOUQtw2+6k9/OpNA
2uOMW2g9ncMEWZjLx1gxJ2JMS2A2iUTZPjrmfo4JTPie1BEN/zxj+umd3vNYn5tdz4VRon2oi6Um
+k/nLccZhiRNqCxN7S6iIKBz6e8VxY8c8H9caSl2rqjq+Of7uUGHOC6L2piuZOaVMCIs3rt0kCeU
rUsZgrlUgk/9JJIBtMvcOIhX68+B4oKX+Vus+RF2blUpFKxUzjoa+sHTMZLnDfm5QbuVKLd1Uvy1
z6n2uo9wgFY690fpHpzSQsp/dJBxMismzaYXFZfgxhrtWOr3GK8wYjnVMmTghZcUvfa78zjMoYjG
6iJsCRasYNdXxHbFHxgDF1Cm6x7+fpZfou1rxAjOk0yxw+0aeEmX6aZWcOCju+gcAFGi+ezHGJSr
3jW9/uQ6pOj8EKpgYYOtWHbmJl8B/QNqFT3cZncVMfiZx73TxLI+hYqlembThjZkNd/rbwD18AFY
7yLYzEVlXLqfH02KaB5hJhfgmWYexUg2AbgQ79LTsz+9a4ITQV8q431Ir0KmZ2g5ApOSI/46kbW1
s2SwSXmeG5MLtlOknwsP5J9ow14KnkcZ8vUR2u5IaIZjPhyXbYE82UA11G1yGXAtL/QC4hHfKMKJ
czJ/pvFseqIu973rQIsO8vuBVNV6/PfBJKkUWHu0Pms1vFFuqYxz7HXytH7ivS/mpzFCfBcedZmu
DTOjrUrl7BotQmnld2JbInH5+K1TxBqYItQ25fdNKLdUFgiq0FjT1NEhBqR/PnzrZGZVOT1znhco
t+Abb5MgZu5z6OT6TEm4rThCIYrgGNLsCAUIs2xI6yhp51cIJ3maXigksJjM3UiZLV04WxNOuEbO
qDEC8F/I2IvMhJ5njs6mCaGWkYT6E9aewRammcNpsA1Ov0FJ0+E5tkl1Ch8KSMmzk2hxesIYknKs
ZAllXGud+XM8T9yaSwf12MS9c/v2S9npuaHoPUUmUCd4ozZs1s00G6bJ2lcpon/pC4oleXm5Wcjx
dydE+HDqs4Jn5M3oWp+9IDL2aDBV8gbpnRue0GChn5bcPv31vi7rhQGSRcA+Hss/odawWQvjAcOi
Cp4Mz6Jd2QX0lZ2Z1Rsd0xf3TYrYtkPj0KxhNLh8RtPmVUJNzRv08n47tvAlEYdM//Er93kOa/Le
ji6nyPNuy1JgTeMmuNKPZmUcFNgobyYRax4E2gjjHb+bWTKrWct/D2FVB/J6lARTPYaqaBMi328h
kfnFpyCjIaE5DVSy1sQdvdyEZagF0S3DxEFIxJv1eCL3710iYPuQSsWqsmW2Q2uRhdxmR6Xq6u/W
1/6DmT5XVS1rp4CBwyHPHBrdwkSOnmTs3AUtPHW6S76OrR0a8sZCMZeBjBHW3jyGHe4UzZjyHVSZ
l92MKm/+I8eRBkYnmqUSngy9eFoVsJJvuf+iklir5VndyHnHHA5f3YoLoJqyAac9ce5JfRunjvs9
kLhsu5k6gCYK44pl9gb3Q2yf57ZEGhWdTIW43pDTBeP6pjq4yPaYd9ZGeeBQajE1CT8eWmmW80WX
SNPAvlwGCgk5UTwtu5TrtBSIbGnV+jqkozthBp+Rm5mg03OPrOI//0GpCSkhvJYsoUibzgk28S0q
13sJ3a359t53bn0XFpUdQYO5tU9ZO6OQsyHR6Z95ubpUAlziSuLEPUCd/Hk9i7NQZKVSe09MR5zb
lg+s07g/J1/SE01ipq7v9rIsK+t+4XuNXl1iLOPgru54AlT5sRILolM/+59e3pT2p0arMPtgxlyT
H4jcsaUUUIOj4yrHe+6oYHt8mQOGgU8xDdho1s7n8hfnMvlNIC9XZq0dL/LGhksjbjy6C8NvaTIu
dxmKsak+jQyD8fCMOHHcB3XqbEJbhYvAfwGjlQQ5X8Bp11b6uitQhg13EeNNXI8JKPWo/WNtJEw7
OFDREVoYJZyMPWFA7m1zxehi08QXOSRuzrIGN1E+VduD6Z695KtZz4uJHFdvH/uqs/0pbB5l2bUK
mKbISeqiJWtlkWap2NpSi3qsP/B1NC96K3Xlu0K8xpVR3RYQZnUxjHCBmTm3wnXpuWBZLZmKimOw
phAA3I9y+1Yp8eREWLMlZDdNlO98H2dHHOGrmiG3TD/zgW/Oqq6gvqUu2P9auHpoE4bXBIOIuGJv
KBRvXjHz1EVhAh30yueoH5NhCJyE5dfjw6WFGHVej6ku4F7x9kaTYezwulV7f5E2+QlQvj9Pai0a
CYOY+MypaoexOmzYVbdjdq2rrFexnBn8Z1nfjbGhXZ4U2TEG4037e7AErLRieHn5nooYwZCu/ZKP
DLcVhU1Ve6bu8rACmaud35B5Qattgea7/FGhcnmks7X7Td6VhtOIDHEJg6O6OS6JMcyVRkrJwDuf
4MNxXpPMv7siroBmx1Dn2KOp1lObAPsMjtTyA3fWdr2q1Yjo3V1uyhRy0xMmkycXmZ+pRSll1MKg
baDeA45VPw2PywfSn0f8+WS33SizXLWs2SNCeD0Ef5iJDYLMNa03w/0KW7y4FYQ2jFFBkrBcU4a1
63g0so52mrweZLEZjqd42AtAhXy9d5MSi7klSt+yUHATGbRJ7XH3R615kjqrggqBuclI2SYAsMr/
iZME8Y/JcjIfrevBHjPmZSH8VvqA6d9pqyF1tS4UXeFmHsPFsQk/phKFyK+i4jxnxuzQvsxpAYTU
LUfwAg8yCSxbpxTCfc5uXRFomwxgfTk2A3uFzokG3K0d5Njt1m4zVCFd6k4fdk6D6n6Ra579m01M
9jSC7xFUj0OWtedSnY9mRRMDFoyzXAKofOoVAD5fT04SRNAiQkDH5hRgw8uxeEuZbpupWgQOW+PG
7CJTC4VHT+bq1gpn9jZRbAVhkhPqzjnaLus5gmAXjiDJU0gk0FmlFeWNhWToPDwI+bPTcsMcgag5
lMB3+P9R/fpeCKYJQ09ga1NcAsjjGUUnxtXFk3i8ZnBdG03yAlANMUi1C3uNTvWdfC9haTg/OMMo
m6P3sCfKeuouwc0yeoSRYhfxyWFjfetg3dW6JD0kwyM1qOfQOWwFGarrm/F0pCfEcf33p32Wd6Up
s/ZFK+YQ98bcLXwIWX2XwLJeZDusQXi3ZeQ08Qygpg6PuCaOkvMEAeMXYI6SdRlb8RMm6LHwQ35h
SeSBgjBqZqnSoA0ygpzRZfMlPH+kDCxfy5I3r9vlVDB4JNcKU3i8SZ88Sycj7FJ2X0egQdtFjSjK
rGmQCtR/4kN1kvokfLb8a7hhUCS7+DNWBXkk2FTgj4mBWhcBp/z3SEMy3v5MQffoPaBfxESvE7P/
qB8knm4hYxMh76Jx7Z1ZIkAJr07UPpyCItJjqvmSFuu+zk99qKPSFb1KX4+kfFsR12LstnBiUd5O
ciEkXBlEIHDKuphNBvuKH/FkwfUeTOZ31ihMdNyGjGTyEyKlY2lFzrbEtGe8RttEsTS56GwIbXdX
ObvE2ue6RHtCO5+jMit06wpY2xD8M6MlIsVUYV1Z07E22++Vr45eUEotfW3yRQDwB50jPni/Kckj
ZKjrabGwuRHCbHrJayO+QhKOd5dAsfBeNQte650xPJyzO2LO6r4xexNTsKp1yLx1YNuBJy2BWbxS
N04xRmqLrpehyvu02l2EX+T+cMHElbaLn/30oswf71y6fJ/n+7060vHXC2CsPmu0W931WzFICjY5
4cLxY8/CBTsLWkulrk6g1a8rfgqfUUXIUhpy02ICdw33wlVMUIvMnpGZiCWQqTevPTnKMkdwaNFQ
yAoEVh0ZSds+DAOEnuiH00mK0EuzxGb3MBOJh9DH52hQEOXNFtv0S48y3mBp+i4jNNFoVhP7JuKf
Tl9S7LDW/q+Ao+QNQxoDiEkvTCgeeRr5Z1v+U6zbO9DDytd4u290n4gUbUZyLcupL4AwlSsBJKqy
MhlNkbCRmGYdpxRqd/K0G7hT495RQGZA7Mfc7ErjRwbKHV6a6SrL4FJboUTtbQ+5/L7FEAJJKMEt
WvxKWX0cM60HD3hTId3TF8mph6nygd7eG9ZFFTvMEQuogL0y8Hr+I+h7o7YjJJaoNIefSQsNxnj8
mbCwkBaiVoyj8Xo/jzdZqbUe6kCFLVocRR6HSGRbnYBjqMySVavAsDluQ+lg6fyZK4u+qcavmVos
gFvjxYZSyVtiggAKOv2vgQBSsoJq0mULoQqLWn+czZDMRvgTP6Gj1o1TnnNzQTWb4k79KHFb856B
2aN/cQf2xIm1O1fT9X36CJSPNugIhjwCm+XuJgVd37ta39lfvUBge8f6CjThoT3oO1SryaDBQmhu
rVVXG7I/C5ZP8q8sH2kxV58rFLyJuxSCzbuOpm0CKrakZmgjwElFrJakmtRFiAWRdz2zvAK0Y4fN
yHhGMUVG/HiRaORFYGz5M73Tr281AAIWSQCO6bS7n2O4fXj8FF++fw0jajTJQZYybOBPnQdpvrI0
yjXJvgz0geirh1Rw59xb+ZbHWu9Ltcusx4WH4TNkXIeHaS22VZhWGE5btkcUAxIKbQMDIKaNHDgd
Y9JrcnZVXkg6MU/Dj3p3ogxGSEBaZLJQXMsZ3teh77v8MbIoEztMfS/0SmuVXoiw4PWvsI4xAt0+
y+LzkDkQLElZqPBrZDfM4U3yy6hXbxITzfB91HOgeVULdNU0AdimfTWuv/cDGdTaXQTKmg/sVnWv
tBC5Rmg0XtdZaqSiEUN/eXFN0PFGVZNeyTOgO8GSmK3GwPXZkpZ6UVUURKCLBRNIb56N09+3C8IF
qAcojdqk+9F7ExhuHBjCWs6xAO1yzVISjrFSA4LCe0olJ/fRxQFItZ/RRUinkQXTidSjf0sDeWM2
38CnSHs5KWILLXejcCYuVRnJelcI1Fe9aS62FN5AhEge2iRho/PYajk+qljlv95XLm6Sk2K9zWGZ
UV5L8g7LUETk0r48VuRVWptO9kdaPRcKIroMTyY4ukDLFvQ/byq/74ccqV/vYDHemetwDwL7TI+P
1/+O+iYDqExAJjVHKEC7hiq4tf5Rqlz/+73CMrMbDh/Jf5xp5YVlAKAYu7OUBFlc+JfnAPxU+6Cs
z/zYFPEPnk6Ku9ha+rq5uQh5hAyr45SCtJfTvwvU4rwIuJaCL00f1KtrwkpFRqkWwPt4gkiHab3L
iE/FuA0Escbkfviui1mVckB4QpCtaCehS6MKTjQUqvgZb530H0VvfyrtvH9oDhZFEkDmAu6WutT2
pepiFtHvluMCtYbUYH0pxB1fIN+Rdy7Yc7VrOw9amxo6k4OLsVDFQoQF/tj2VNp8L1h9JSf56nXf
0EDmQlQ+smfE9swiOoTbdPpXaq20q5Th0bKaVJKHQItBGJMawLDeer8I0USnmlvcvUv/LXlKJl8e
2k6n02/bY6B2xI4QBrRVHugEU87lHOb8tHf9w65Pcttc/tjY4I2eJAElLDMWwTUZud2Iek2qy+Ao
Ct4ejSwmKzh7/dljr5CNf7yhLomErJv4r7GE5HFZhPwvkaYlHlNL5mgsUJ6bJzOwzfILYHbwVl4X
rGV0cr7x5S9UiYoLLpt0eZ8EwA6SPAeqXrRHx1+hVFm3v2ZcW+ib/nf2sP3As025HzxYcnq/WUGA
qeWQ2zkx9eTad306kWtMk5fvEqIk/VxaEuos9M+ikDTpxPbnyBSJlXXHCWsYK6D3DMtO4Q6cSwDh
/ZDr4BYLHKacfko1jBj76U6eX1NiUsprmFevMHC72zAyG8aI1iIx7snZCwy/H4SsiUISeh/3CsTd
ooNcdiTU3jKC+lEwjEazf2krck89bCc9B8a0Hr8jR9cOT/Vv6QMZhZSHuY27ILDNcr/SBCY/aj27
3a16g9oE7Cp19LmpTbrm/T/0oKBhB6TGP52/z6U8umst6IHZ8aBAYrjv8yzVwlcFn2T+qgSi1Kkm
cIOriw/kAvsVrrjOY69oih8DWVa3bwitB3y7ch5rfeqTLkpEE5qV0QHDXnGn8SZXxzX8CKylInf2
qIYSRFmJQid/CtKSBEP89cqz9Eun3fEoAZnTtH3vTlJRcTGX7V2JoNuvQlhcfrxhRN0fLh2xhZTo
tgI9JrJm2WwKez0gJ3MT/gIFARhG7YALXy5YGfXoObDB5yOJeHRJuKBgFOminfJpUZGTfVx1U4V/
iILEN5wdJ+MCEY89rXsNgOxfJsatg+r+zpTKZKxqzgLF5NWBXjsMMnZkAWwj/BweDP+Mk4roOLlo
JVa1mGyY1vQZ9CwYn4lJ5eRi+2RkaN5EHEHl/lSC3FzKkrxjSZ+UFRaBO1v6sNjyCHUN6Z1qamdd
OGmh18Z/DDQ+WqEHJDZS74csgoHKUk465baS9Sgiz0AXBzBMx4eBUnBfQUBzX9l6MxG+l217zgep
JdLkAtAxJRvX/hnFlh3Gw6XgkFm4za14R4p08mIdsNjPkCxC8+NKESXH5U0KkvkkfP4qu/yrDR/l
CiKnFFfBiLRv1nmc/mZGU7FQJjyvlKabwCeCfrh4yg3/01AKzHB+t9BLnRunrWWqPNqXUAr83gng
opshYTb+WAL+38heZ9OpS+BuQt+ASYjaZf2Sbq17wwfr9Whb0sBGdScFO/4inm2iU7gJE5NA3oez
H+zJcdDFNyW2mhxMxMe5A/RusOTgGq3qLzh+bOK5FkBzXQ0Nt5XQAugdXUd5EvQQmzzN0uD/NfD6
K3xqeg3Fp9XvCIcsA7nQgFqOZleRZuDR/4cZBaumDeCRluFVDtL8Vihz/6IZ5+ee252XOB2DebKN
DK0AiUKZYiky+dzLeirnmq462s3bLJhfDUiWAsoEksMDKyepvcMLqpjSWvZ33wMhaS6KeWpP/N7N
bmSaToqDlWHb0AVc2ozDkH/H9i+IshHyYc1+LO5puM3fhA3E9YJfdgcZmMFALBz241KpMq1vEUsN
+CBITPh7aGv494GbquMHtOJDyaNrybt2FU52V49XxsSwNIvEQL9gNpXDksSplj9EvmSpP08YXTfZ
YOccFQt2Ojnp2ly9+KnZ5MWKEhwPp3rTxNG4/Pe8qNsJT16UNDjHlC85qpHfyvK8IqN6RGcQPA+B
6hE7K/0Cqx98K0qUgnqUfMiOKbe7QY01ytgFCx28gAu10TZ9UL8WZNz3wQ98hjoKXJ327wlgP3me
s9h5vzgPCRsDiSx3PbeZ2MeH6ks/PHSsaVgDCAkQW7f2AgC6gJCSxaSUtf+Fh7I/cMkq3Gg/yCWT
KNYLqMbQgLfo4cQhmu6Ssf7QZJ6F7Kpysi6y7xve6a+SOkMc4rgnRFNe+GoZ5nj3l2NKMibtsKRi
d+N+4IGIs0ersxs+N/PfL3KlaeURlc7MO5vzYe3OGQZPJOwp4oV1ME5sy4sTwLE4e1y0+vDSP/rS
qDiWKMSpESO+3yNMr7TyUawYD8BzrjXJKSbCIkwzdCeyOh0bOabo80KQazNFqIQlA5JD0QzeNiqA
inpqioCV3WmQvPEBh5zV0HaQTYFfZPryVtyauPc+Qpc+BsEn69KSRUjBjoVItcTxUMdcFlZnMtjK
4j5VoFvCfWkJqmILkaBt8yp33nW3mqgZkRzXALwWBP5rhdV+ZuebsfszMEBtLfSqMKoKRVmaihMo
q3SZIwuDFA/egn9Sgp2tk0G0vEsfufVWm4CF8xXP4JcMxfmQ7Fp2kRgtuZpSbGg9CBdrSpE7tAjJ
dTsrWsLYYesQA9wEDY5Ted99REaFusqUJu+FT+NG/kOSuqgoRhH3iRrp04iDPI1idaKopyt6//06
DZtKGylLxKWSlPGb5FPelXwMpNrHUW//5Q1Obb0URv3Vj/4fGuc9vTeumlNC3S924+oWI+P9v2PG
RYQutKJOWN0mzr0N8yuHUThN6q14QyF+3ELdi6+vpP6QOugRWWOv8gZdhglV3tzI+MkvrVLuZ3R5
i+BiAwr4pK19hm9uloF46TEnrM01kUPd6Tx2BxwZ6rVQQG3TxE6pSSRCTGRjP/Li6p+IETl35AXI
p9XG/fSYC0eqROZ8f0NXj4mxM1RizRBzx3ZFO+Mu+S+R0NJSWJi0w15+mMuoCesDaAcnbG1D6nuZ
391mOSIAtBEkat8ITFYGBN9vuIBkdSoFFditgYZTCRaLJiAB2t54EMuJbe7d7Pq58krXaIVAfaoF
NGMZNmD5+rf93F26VZ8WsblV5E8tFUsp0ghr0RB9YilDUIvBZttnjxT4mIkuwI6EVaDxmSE8ZiiS
4pLyjHLdC1q4d0XwpATToVUkaJU0ib7O4It13tNHWaHmlHLJcqzXocxTYbjr0IrC2huX+3/+1pJZ
aLhASLOVEjsKVHKdqxDw66oaGrpGknyQ3Z3ifbMQDUeECXXu0+Hl9uN3kAK5qIBFhCcsjEput0xJ
Z9vQhloNlIRRZfxcbhuucJecv33HEoU9KmEUcs28T3dwPtSbjE5S5rGmIFmFXMD+tkvmAuUMan4a
gulsuVbkgKI0dOSj6Wepp1WbLh+SDoNJ9GemrHA8wkUBlZOwOxb+bsOQHxBscAwu5Sa4i+EHowym
vX6HAOxjxuxP6wNDrCp0AbyHD1+l9NGlNONICojgpHpPBB0kx1p7wWEtolpkOUa8euW0ZKyqzvEd
qjXcrCbw8Q3VEkUwbNfxLibF805wHnYGqrdTgYWieBJxadCcKZuC6n23EFvzmkKWBIw6kVrXascW
bwG6Hf4frwwUEclnBDBHC1PJzI5iBiNeY0ahCQswLXLj/bpwzz5E0CmtumIyFlWX4P2N6FYjDd9I
DWcCUSM0hDQepKHmBChs2y/Zarpc+OY3AOBFDL2mTdgA1biNXk+gcDekUrkEHG0q/9X1J/oR9svH
IarBqNRU/zQVsx5pRTMNyElP500rY8nDgrGAnyLcHxh0Ra4i6V22Jmt/o0XS16R61ZOxscXMfU+K
9RHplHqkeyGg2E5gnfMSnJH8DAMNPeAduQBgRdAjhAJc7PfFTjBoTB865oHm3wuEXYdzlRFAjAEI
Bqbx3ERW+6PM63TbY/ofn9XL1VNA+FgvAml3BD30Ug2mHTexxHQ24Y5JGljySmTTuQFMMZC4xfHx
HGDXzUaSQJy7BiMWUJwANdy/Ox7iiQCiBIGbMOoAqIXdooI1bh+Z5oHuSqIyNXHnw1WiFUe+OFif
+K87Emu/5sPuYZiSFR2TMTK2/ZVmSvIGtWY9vfDQ+mrG4gi6v79N23D1y732l8ICJpBe5GIPVLp6
bT/RACwcgBLYqwJHNWXLfayhnj2U0/fDiRjBM8MrE0J24hSFFFguiqwDJDlloYE5RzaStCNhuA+o
yKAlgYFiQT9cJeYdla/+QeDM8C9Mo6MbOtHyyjHgzPJgeM4jjiMWKg9Mnal2KBy/A9CoEIe2gmVX
nkVeh4gCjNSsgpVlypsFZ87zf35AShxQXn4p25M3uZT47mqvYzGOJkzwcXUzH9WIpQdW+99uBzO7
jZqJfEPyOVM1eZfjk3RhglOMscPfQJSR7Hu0mnnVPFn653Da7OaC1f2amcYyf6ChhCV/NZDoiD2C
xQg/N+PMuFhSZFRkVSqqqOZxhokV9idGkCUJ88y5eJbG/36gWW+53aQ4nRmA47RQT9sN2ipAy5js
NiGbn80wXKHvqOeGIKQM2LMOpwHq67eB5xfO2/5mm1QVDuMmkakMoP9Y0UKyuFuzfndgJwgecLJr
ebWdTZpDOsrTPF3UO5sOPmRMOq84qT9pheVoyHV81+DAC8O+TR+5oNxa4gG7XO4deNo38FDHvGVy
kGF42FvQHbAs6dOCice0ZAU/J8C+NdVJv/Ymd71d5jkaAKYPMSPwm8FT/50CaRTr7UT0DWIRV1V0
/k9ebO5wzCrEqlOT95DhRWP+SIVip3kViBgLH5CX2kMeJWCCQ56N4zK9rYrJmUK3ZKVTlOnrx5yb
CLeioCxz4dO/tN1DuU1y+HBO8xgZNCltVqc4mMFhr7CGfsnAlEbfWeh1P4a+KGrLmtdVrEqPk1cc
5hZR0aHIvZ5eqPy55PyuRxH52Cu6+52uni+BKUh8n0ddqImFET81pYyDRQhnLa8fVRc9d/9tUVDX
bh/YE6cXEOsjHLVY6DsG0f/6f9JXfo3P2z//HpiH28GYtxm2t0fJ407exWTRm1GxgL7dIN+rTqpf
wg22zqBDaS/hFrg3JWTKoG0Rcy8mPR3NF486qAhtNnj2Abi4qJ0t8H+eAQXJUAWQzWqQQ+pbBf4H
AFHRKx1c0i9AnEftSY/HhxilEZxgWMTlYWNSSYWd1ueJybD+TQGYTUH8Ap32NhLJhqNqYY9UReDY
e5JR4+hgVivbD1Bgj0ZGjYJAL/vAofY4jT5AFFE+ZcrGw417cn+0b1lF4/gUb/6zmPOst8YLFpOW
MHGidhGhnSJHsX54GSvg2W6qWiVMbZLKwk6a7tX7c3M5LaaWtlF6lCIH3rmgl+YWuuxsgz39bHdP
52yEIncrCQ0NapJwHKZt7V7SRqkl2hR9PVlC2je7LSAOw9M6n284N6nOlFbwhFIqSJrN1Ukbu5wX
FQHQeb1/s0JbVZlCG5Cy8DMxXQyRhUP8IeS51fL1WATSBn7qRUv7Y693v5XoXWm/7591rL90Ap0e
ZCDsB83ESlYQJUWTnq2mdkqLQ7twiAHLtQRAsK8BPa3aZWVo30olEKp8TL9strhXL6YS5JxXjd4K
htLXM+Ypv36jAjTBGxLzuzl5nHL+N/YnGJ7435p0bMvuQ/d55uwWY9xQZGAV6O4JKtEiV2QLlyAy
UpOoawRJB2tq5el2ex6mI5uJC2IL0UNX+/JWOSNLnREv6JZY2pqlspWllnRPoMNQbhEAuEZjTCg4
vApJzwJLUEKaxWJycJpzhdFBp7E65pt42BkZCrhthaTmzFkoJD4/IiIT7XYA/Wnl/hC1bOJGGksM
Olyh0FgSmD8nhUl8PGuB2WDF8lsbwjRYRJY2hnAd4JuQLf07C0wsnFVQMnlFXBm5H+0nry4VyPay
5Lgrlv+fKhVTBgF0s2XI7GwkBneOZ1j2MdbyvljO/mrmu95mB3H5JIBQAh91+RhwkMraXP1aJXCS
K/6ehCdHc4yyvFjLHlT3WMB05Hxn02UD+9xkajmxaa/DIsA00B/LSzNUoyKImsPuIOdNNOjTVyIO
0qJxpsNqbnaSwIFn3DrUEIm2mM2tGw5yfTBkt+xAt0DQoaDeCTcqweaARC6Z+Rg2c+HczS6o8w3X
Nal8qPU7A1adjYw+mPNK1Rd9W1RmyljNFaKTEjkR0whvGmRAOTsYpQB4Np3zb50OSNEBcZgM4K17
vfePTGzogHuUyAZaXa6LXrLw7kUKowZuja6mDi2uXuRIzs4potMTFhaBvxranfcnJHp2SfNtXaSL
VjiuisQzzSbF08183c4GwB7II6tjah7ifcEEjW/fC3DE8VWynW4zaAk+GU8gmX5/CykLYlLksnW/
8RaJ66fgOm5/lK9e1pLWfVERrhgBmPzpzRvIwVHQwUoZ03xS7c6xg8+4+OON+Z0TxIt5HDy5wRWs
NTVKkeFSrPSLHXT41z9V8YGfZEpe7S6EdrDhfFlFyv7oT5z51ulufDxopGDiA8Yk9Ya5L4xLhkA7
sgeeT3qHW6wHnpGpJOFBNicqqM4qfsmuIj37/jD7T/7givAucSaIVmVWUQVAlFJPfvhMa8tEhQ+E
PiG/0xqFKQmNJBlp9Yqx1UgytD3mUTB6/XitUexlhrSwMzeYtaPSNdoFng6K8ljB4kvx+OMhueaR
XC4JwA72oaR+G1X1UPj+B4q8fOBK76E+4Zcq0QV/k1PhJtYYpV5qefq6ZtmAskGjRaW/73jO415o
E7pP8xM9lzgN8Yhr6bHLOAAnKWqQYCQPPxBGVTpgIAdcf2KZ7gGaxuMBX4AIOkli+Vrq0sjoN5wp
B/ZYyoQUjEuhD9YYT/ZXRE5Q79N0S3XuLH7u7yKkgmdYDw7PqjGX9wQsZ1Fa21E5fzDYMgIlYrPP
MBHB+k5a2YyokYLfeq6rM2Pdr3UAhotWP5p/biHESCMm+FJiGxOAdFrYS6iItHPYk8JkKJDUFyhs
6TB54aVpHTq+6N1aBv5n1H9rWkD8y3LwVRy5KA+au+EQf8Y1q/DOiNDLAoNDon12XXyQx0VH8Dyo
bad1hw+X7mkLetdK+PYE/L3Q6hYZCebZy4MDUVNJ8ueLNcYkTVoqBPRAkATO2ZPj/XQXA/Au1gWi
cqM7oCmCwNOPRRG/YowILSUFh8wTYN11Hy+oHf27tHVqFZmaN0Lfm5sO6Ingk681HkyCkLe9sadz
c5USniLuTYP457s4wPtpjet0ZIG26zCHIxhwQasvaQhXPDIV9lKNipcjcJHl603FZ+NwNqtnbf1J
hnEmNmLBkK7PMGlA582PImD8hOsWnglmlHFB6SGmoH55lJemaQSu0QwB6dnNYcG9Rka7eV8gdYdc
pW/jBuBUcR5axZJrGF9uYJ+DdtpVnlKIbe927oVqMLohEmOieyX+E3OszIzbrtC4udec1FF5PMWm
oyDbXUkFUBd63hDW7HSxJrCtjJj75xLLDAencd13NW2n7H7Iv+E/+LYAPp28m2BXZXlpQzeu9YZ6
w7qeW2I3kE3m1We0rAPZg6JTx3nfz43FHlytx5x/L3SL5Ur9oHR7LU/KrtqGETDaqtshJ2G1hfA2
vZV45dBTM6wkPE2WCylFVuK9zjfM/ePJitIqostXmTuwxUNlnPGAa9ia+lXxjYgirep/x1Mbp8IL
fZmNG4Njkk+CZuOZgqX68WyDoxNHZXHa67Zi+JoY2pP7aVvHZa9K1g4jqvnULg4oq3GIUx76PuRr
o+R6ikJGXqgtopxyaiFYUdpsuUBGs73mm46B3SWNLPvSwjsYIpa/rn4ywwXyGVHRVUco9BQVNoHn
HDJu5sWk9sDOp7tDRayafCZxovkRr5By606J30xknryP7BfaniwYAMAQX6PI+8faP2AEeXvuIVo4
o+x4Pbaduvqxp6JrESArA1io36+1wDw6rxX20w6XaST8gQpGhGSMStxFKOfaIYInfduD/ZlbXZrr
/8cj12yKSjlEaaMgpULOc9VZQNE1ykFvpw3ZS10XODaTyWLv4TeV5XBfwlNJw5Qdi4AwktGbDo9q
TQqy5sc8nSxHE0Q5XBntDyFQQVUDugt0a8zPHcDz2dKMxmhx81RI3hZRUYbxc+zYT88ZEQhhe62m
V123RvUmOqBQAzfcprGQO/qDHzI06GP1einJJyqFh4XHdTYDdqCGZyM/fml0j6ThBeggVA/J3YbL
O3oe4vbSen4e3UsxfICP6wjacIMNFuKKcy9+a7GOEnwOwKPOvL7TGpXWWJYoWCgzxJ4A9i9clCPZ
XTD2EwWCZsoxHAw3skMQ2uSHepA9BL7S/Lryi7auNkzJjJoOqM4+orZAKASP/jUOaSFhoegzKmxG
jSzSPHa1bYfcCuI9SDycUDFdEQHCE/pOAhIVRsINZ9Q8YPdVtInymUDy2flDgXu4IqLYsboaIC2c
XOsN0GE+30r4vDZ0w6yiM8efKWcjptfcbPtEq5Uby6FIkFsDl56xPOq7TM9nRHI9Hdkny/69+baE
76CDXRvgetDN/JhtZuvqDbDi/sS2r7d65G5G/mPBPDu+u2OHip8y6xEbWnmBi8s89pfqzzmJrz47
F4duPcbpEoQchj1pmjLJUDqlySgDG3/pvN8xUnG+STrcJXkfrX2zPRj6PvQTBIMEsoFJOkYG7b26
sTbcIawaUuR9IcacEh8X058CBwyf5U+zNfg2xoS6mfbvLFYtQDFjn89iw4zNpI5mZhc9XpBt1N8H
QYD9gvyDnfTFV8w78WZOcSohvlb5K8DlglGtMLGAzaaZ/IIcIHl0C5tj+ZQtNlUuPrhK+lSHOuDV
oYnan3AizsQDEo4Kgt6yEalBy4uBP9I4gLK2K42KG0XxaIeuRyMIrq4K+6gtnV8/vwnDooC9DA6G
Thcn/wA/MXz6Y5fMD3FLz3SlifUEKJyIGr/jcpBM9qnf2zHWQTuitrcc+c7H/2/lnj/na8NPRAk4
kcN7G+D8CtIQC4FT6QZ7MnL1yHpej4zTMWlO+m/7IbrbF/zxDgKAkWSMZP9e4D8Y/xOktymj7RCw
I/q1tCWFbtAMRaFEhDbcfeRKLmWw4AjYLsvSvc3mV6FuLbeAq4HA34DuH9hU8iTB0k5HEyCQaM/z
qAG9KcYxk0YbPX5uiw6ROADMR6NoVkH++l1ymzmahUGRAogxLxIv/exOkSEaNurnVbl5+Dpbqv3J
bkuOEGzLS5Z4SOv/Hdiz1d2ycrCvhLroli6wFIcZzWZ2mlYDkhyjtzT7kmodAofISHL0n+KXm4cZ
zohKvix41BuKcMcdg059mf/BL5Oj7pI2VkbASfwzGfTrTRrB1B1/HXlclza3svlRLm+XNSUu8Yxp
CAi3s8WD47tUeCetqd0XF6Ms7EcDYJ0dF4eP4uR3LG7EMO5D0+7PaBv+U3g8a+zzEpC5jJbted7o
VYbvtMHrQa3bXIgk9iWd01wv1AuvqLR9eVghGql5eqpt4qJ+H663ili76Ao1g1/SPURV7vHLcNxr
/zeHx5xtKZxslFeY1N8xPzuTYt4N8D1JDEWBc7zfzzP1Iqbjz++qOyoYcfoSpzeqLnGzOyC3eI0p
MceECj6bqTl3gpahFqsWgnnZMkXLWx4GbHkjhcI9sFLmzJr28sIP7b/A8qKiJBF0owqDcBR2lINg
elMG/fgyL9cjgWSuZC2w76c1/C05sPPJeHfEC5talslF4i0LR5D+e4W5BYJVOp01Auoz955bACvH
0MMmUL//U38apqXIztpX/EMa+ES6rfjaP5oQym6ZvqWTEkWX5SZGOLZUVJTbC9pFkkx2B4JoXCyZ
8+m6rv+Wxoa/rEoSU3oPiJG6TfWXPvVrTFwSxMgKb9ZUawHaV5HMZ5OBe/BkP3jG6r2S10TPYWQp
fRgpFRrY+hXj8rbD/X/AxE87szsoy5PGiMukJRmK1lbdvHQzZ7aziGDbiI6TQGXyi3fMzXOH0elH
R7Hti5fA7h8qJ+5QfS610eY72/gSxPsUniJHDqhgELRN/sfOM8OG2fHMMVnMtcEQwBpEk33S85U0
iWcYwk3VE/JKmslRhZBWJnk1B4fltVmLWbL/HO4xBEQYCVbnd5hXtIIp8uSHPNh3gprzlC33G3kC
tholDOEIlO9Rtd870T5QnqYpQaWV40QYh/qjyyCVL6daxG6uhS8i5uGwxcyayEl5MyWBZ/yMYdGp
hoEid4mdplXVk3hFcSKI1GGbSCqLKkujSyJCjniaJatW28s8z1qws5vb9h5n2k06URsJwqXSKSBW
XIr+7QpclQ79TsXZ40uZyYQvyGQm7DTBf5EowwejVq0oztUs/K4TMH7z1vzvLZW6qyPe9YcrtGXL
MKTPTtBBhz5o09dZOOYC5ioD5OHLA8h45H/9FokjYMB1NaEaooCiu18ygGlJc/LaEnkx/UPN3FO/
Kd2osYdVVFGV6zm+uRPUGgccwtGkVltFbKmO9+dvoc9jjX8Y7cqhUI9pAnP/SXox+FRX4uN1B4V3
lJCo0bl1LI9XjCjo5xaJLPh+dI1x8duuP9JAHGQDxu7poIBQzq9qCuczPdWAOsMxXHjFGaKQmTRt
J5qaWCrIJAHYkSr/9iVzTzaWpdrj7e9P4RCa2xdcZpD10f7JzuF2ZNMXcmAUTt9HCdLiUSAtzQ1S
YLVn3V13GNfIJ/HwWAy/zKXFBjmBkD9a5UUNCD3IOT4FVUs02EhfhXl9Xrzxb+sn74GNG3uyud3U
AwB6Z0nZJ7VmTSV2CP4UzA6KADq6v/DHpVJy5KE6Bb9V6WD6UnmuvPT5ht/JF7kghRjyDGi+2Yt8
0tTOXC/xYZ5yvehcar3qA06PBitSsoDvxcp7xJIjjngBvqQbjHcjAFtLs/kc2A+lZLHWOmRGOKPg
YRpvOt4s4T9NZtdu3jWChpMewm9bKrjjzM7XkrbL94baUROb8SN//cylKsx89JHqgJlOzuR7EXoN
kJ3CUMojazBtA3TTd+5VYnx+2lMUhQnXCcDUNlk+m+kEcX2jKv1EfHZrPko31ZCwXN4x1FGfhiHw
a83iu0lPiicG3HJmRb9x71nXeLZsk4Rx6ltdhP6CyEOhyV5pBOhCprJGxwC3h408ns0TL4viDfEH
ICyTmKWUepVInJ60ZFUor9FEEQMPZYSr65aBDDhQkwRYht4VDHqAaNQfK9onZixrh1g0ZqeLfs7y
t2a9UJsDbUW/Uk/8Apjus5zcdsPCbQeVw5q/pOKmJEcuFZDrlvPJ5jS/mpqA+P1UQRDJadf7q/qk
RScNSyo7XcpBwmBJEpCcmgyxf+9ZfA0mq2zaQaRLGV9Tw66RCdgVWJqWtX/G1xctEI5Wj8D4XPIm
RZEGwuMxmfIfJIUnOlL0HL+wN2Pzlndgymcit3YLBk8LLIHc4QtKcamtXRWPvxfLA2guY00tUgh/
mHyFVjEZIPK0qohFvxGDVQj1ec+VQOeHusxDDlSR9goHQtTTgR19b/poKf50e2lKweLSHLLXlcFu
PTPVyAeUpeIE/kx16wOADSvI8fQsMxYA/ZOBj4JQdLoTd7JrqkvB7057FcGkXFcJsDYPHc2pxvG8
9I0/rGiSCNChsj50H8xBE4F6tEGr4pg/g6sihBunqiKJUCeF4ABORYZDhyZ8oIEz8cKqp+/qccmi
/JM6E1Rhqhd58OVXHgMCqsqUZYL3xn3wT4lperwC9VivRyVrBWwYa6p5xfpgSIyt/Q5kVS+H319p
uyXSQyzOMurMs74d1kIxrQqC7vyIxnCWzhE1zhT5DwoXiTSdkti4UIjv/QipF7RcyOiVPkqRsLH6
537Y3B49lKDIVNVwVI/hrFIQOZUBJpXlLTMie7dfj5XC7KfCDIegoP06yam+cf+Pt8WOV33Ca1on
AJUEFrYpdtriGcJjx8U8t+KHP/2Kz3TNVacTCz13xVS9OXLN5yzgKnpYQZTAUQhPPMDYqk3maFa1
DB/jAcRXEzHl3HCszSyekhniCGMTLI6lt+KtzSi8k9znEAVrL5uhOlN3eGL4JW8RNTnJDpo4zAYq
fqNn+XhmaHtQ87IdqrcnlW7tlNPF6miDda0mknN5qEVV+U+zlESsTtKLXek32c/Tav57akZvosqT
wbNmMBFegfMZuocq3185cg7IU538XbtKGhVU+IA6XTSD3SNoEsuumP0kK/eVFvgdn8NQOCc4Oy38
5mIC0w+i21R/30PgFV9vJuw+RV3TG/lbx8HBAbhjl80iFOZt/ybywSMhHn1ZvVK8vouR5kMKMZvf
VLlBpqvMAiCANAihwV/meIXcK6MnOEQ1alh8oBiZGsYWwU7buOsuObDEgP/YBZEwPDG4QN0JHklm
9FXAEBiyUnt5IQGUSZTTRiTrNQQktaOTFDxDrSgndYUZAAoj5h6rX5ooSewt3z8i5C7YsntxPZBR
N1G8EhB805PnMdnfvqn0qVXao/2bCRn4DuIv9xeLDLUvkqBIPddjUlJkxoZJheNp8C7L7nWdbqFE
uk5s+UgFOmuHqKOyKLvzsHkhb+SU8s9QTQzV9XpO0GTw2E1pAh4+x7OZptJ9CNrrDlVWvM2bdZ4K
4ekUUpv4GzJ87A7sOvWYlj2sXmNDJ8xGVc6Ua0VpCYhqkW09fK0SexdggtLp3SStwEsxr22GmAxY
0OQvSC0ocp4aJ+2X6BBK2KDcNZe3EnGKaO/jl3yMvkAynwg4rtGihsexKhrjFfUxY2xPkuFqor16
zdiun+Mm+yxKC+/Zt6KM5v86ioK37Wr0ClT632BeeWY9+X9YgoGrNsvaTK2OJUT2GJfPMGO3GxA8
ZZ11Vbgv6NAhH8IPxnqW+hSIScLpzG3dVQD8LTMtAy7jUbezPOY8eZ3wbCjUDg4jGzA3msvz+4gM
MK+HJyO4gxi+bsQ3N6+A7BNLHP4vZeA7ljub4SiCB/aReIHGhqe4lCUCKIeadbiNc7T67TAH/kID
fK8g6wkXMkmpdOX0XaT6thXqOD9hLWvAoH9GXVgivSBIAufHxWgNAimEdbvLscn+Z8nT2njvXuiA
qUMf+LRUnB/FlD7tX95C4IDyfvWCBkAlkWKiTHPNsp7o79P4TWh565n1GPimkSBkbIH6QQCyxaRt
WQ64ZiH2G6l9akQ/DeO/nMXMcr8L91YvpRvpIa/PmnYiOoy0bNQ2Lc2yrXuqcf1LUojAII6EXbw1
CHcgleWLUafGBdkYnpKWz7il73ThvKoRhf6lUUOlrt7/T4qg5ERhVXs6KS70Hh2fe1pQnTBLFPOa
2jduRqI5HhC2tZLdI1uP1JexHxF+X9qWJ1LCGT7f6XJX/hAP9XcxRencprX7VP0stZNnJ8j7H45l
qLZQYmR1PC/GP/Yet86HGci+bXwt0jxMOTx8ehBW6PrL/ZNFumPQqp8jw1plz9Ax944+fRvRsLob
XiZGMxoYvbHls8qOWML6ixQu0SjL8jFdXlzg+rfQgQL18R5NSnxOAlzzLnJc2BTcT7eoHUPgSEqK
Q3grbwrGEqn4DMlHn1PNjKvU+gcomhr6Y0S4QesF18fOOlylWx1kH3fTrhLWxqDf39T9l6mbXXzc
bHvUjiO5Eb5AVv60DU6pdu+bfzTtoWLMyoKroyV1EodFJ5nuq6HgnY4jKgp0tJASqPHmnGhbwUJ7
MD2djl3wbfhsfJ/k9dlo2bwTHlLE6F6t/CjkkSn9lYCVl4DEGTB1oYqNIB+iPeK34E+pSxRCX36L
0HT/b4iNZhxWSLUf4RLzfIZbFOmPHl5kMzNWIc0VVj4G28BJdISYbhcp+cLdscI8UQ1ZHMYh2i3f
ogjTM7V28b+ZYW/P002l8vL85FW05KH5dADL/pkpel0RvW5iharZ2FWxA4T9X/Yole46M5S5r06j
FQ5trJ4QPKJkirDs/v9JnE52THiq55nbEAxBs6EDcKTD1FmMoycFwv98MGupjgB4nNGIOiHblaFi
7v3TGzOr4Q7wgpnkpXrx3tUONuMz9mM8CAs7pdz5LhBnVRqLG4usGazmjqVSFGf6St2pV0jO139D
AT7mdS2lWL7iPH82AK2per97/AN8qWfCRIfbvD1X5TcexJEjcMrgejgFDPe0V2q5tvluxaTQ1MTv
RsggU0cPsFFWKJfu3NZY0lvS/PMjEZPaqOrg/XW7jMpHOXQOQ/BKPGphbUdzJFoCxOxpDfj/8oRr
YvtwELabJVvy6JdSYoxGhc1L9nAVn/R+zkjXzB1Cymr0hTCx/NFWBDBT5TZT8Y9ftb+jlKXVZPM1
Lq0/Eb/SjfB+upeQSyBrreeSC4F+WNZF0dzZavwmFr0NUuwFsSwF8/pP40M6rpPG/sN0Ggp15Wau
/Z7PnklX93023PpnSU+6hILzN85yhXOLeNfw+Piu4xY7/aFEp7wvCh2qvVMH+DvUj05s7yGRWB6D
UjOh/Ga58qR49yy3dJUSryaeqW5jzC3pOoyeHF7upY9KBwDTp48a9DUZ6+08Y8IDkmW6DNc4S8A4
426eljLzhU0w1t2z//QjFTwP6if4jsI8YL+XfjOAAelNCfGv9AeJ0TezRtTF7mcG3Xo0GUq9xr+O
v3qBdROuynPd1Bav6uK+QdLl2SDDqE86okuS0VQZwWfF8JvaOGxhD+ztSh6QMYhzoNS/W5ivrlrz
GGr/dnErIYsAwYIX8Pfn9Z7/C7NjN8GT2qU5/3jZSnlHbQTR4KueRkd0Oy8ArWxqhR041x6AD0RS
+aOwzkQZmDIneRtSSB5SKp4h6xTPKzoZYOZvEb7xqBCfqioiwcAi0NDcaC+hPRUd7yodhhbjuYIM
9Bo8nVxjh3P5hGlOkFfyJ2/NVX1GFrvb6qwsFAHeadfermlYxy1KucYW1F715oOwIrB4HCLtksiA
u1T2ewGVH59SzOz8k//Jv/7Xiu8rAwS8fOb+PcUaTKKC2QzdT1l9ebGROeTEujMhwm+OIk1wd94I
+uzZ8234KdPcrCiQY8I+lmOUER1SWtQz4Hn+k/lrUXN2Xcz/1XiqiezxhX587+7DyEynbYheN9k3
1Z7Kf6CKxOa0sEu9sjn4vTYqPLEWDtv//7lTn6+EcsJhllSpuC+Rz2hpcqWOGr+fVP8iHOSqhBED
dtePgF4hB6KoP4iCivCSiKRUMq73E+sKV/f+r1pu2vXQ0hU7bXRDSsTp+ZQ10PhYAKHjPafhJh2O
p4vwkt0Uh56VJqz8uE7EiHI20cCTYp7KmR0dLenKneijb9r1KUllNHEADWS5yiC8of5zETVLh07W
fVIDTffiVfrHW2AtjkouCtgGKlWscdmZJrdEZhyzItMn1oURwLU/ViiC3PgId4uJVWvSlqTAkDms
VySjG3y5aIdcuTPJJ8twiLIAS9ZcnklX+D9aoSRZBm/2kg5y5Q2ikO+1pZqJa+gt4hYG66jTkENm
hIs4gYTKwiQSMVp3PuyT8ZAytsYEzcWe6YGzMr/tgN8VkDOdiyJECyzUbV78yjBJZb62dqxShBc5
EGYZfR2Ij5VaFDQOZ4O96xKtwn/Df5+hdycogH/VIqdeMpayRJkEhByZolNQykgrHLb1Tgx3+rq6
vfmM1ZE5Mai3IVk6idzPFNpmWrepThL02Oro2OEAT3b5Wntlte54cSY6NhC2wIoMpMV8j9lv/Lis
UzqJxIUussOWk8TyL4XKiWyirrGcemTqWAIWl9tUQUv2VTSppJ5csbHDQ0ido9IS/RjONhLhKlxk
R7J06XycM8y77i+JC/XhhnBowdq3cQgzDfNwoBD5dh7cazqVa8RsGPkCtksD0axZ8qfp+OzMAlWW
LuRbjZmr2AsRuC9Czmeehei+xc09egncds0LilLaHhpQ0xzNuSHytkKn3uEmrTk2BCrzYv0VBOSk
6g3eFzWAlN6BsNNwrl5W/eKN8W4V0CzZrjuMA8ntYLQnhA4I3uZ2zBIkb9ER+1odgGLl9VNKQRma
L5i2qpg3tVQ89HO/DDpl53wr3zrO229O23zvOelRscw8uusLg8C3Po1pab+LWkQJzhatIS+KJPNE
7PbbGwhRNqXuQbi7Ay4SsCdliRdWxqSfhACojHd9c9idk2QrfzU9alcQFjlfGvEnIBbyiLpq72ZZ
ruV7BQufG6MfNfey6/DrFK7d2tAOKeVzsb0k3ohZg11d6Cgsqqhg1SmkuyDl2NoeecLTDtK1Iz40
RgcwNiFQuLAEe7DleYJGghdewcO/8+haVs/dWPQCO1JG57ul8laPZf8Qu/nFAjx8O4Z/KU1DdfgO
67G0YdQ5ZFVyv0r6hdzwnqY5jWN/sA/wrOqrgGwRbwO7Smu5dPy3GzsgQ9EdSOSSHGUTRJ9MvxAe
6fF9P8fzv6nmpkwE7nMiNccpPpy2OGqyNwsVZFmHhA9aoHaBsHau1C2yI3+Sl895Cuqal3fNoPr8
iS8FZ4/C7UkjoA1Jec0u2srXSRrAey9fwejIYrCZUrKthUreFTA3fkCd9TUV61HAXUM+DJPjACpW
0vU8ekK4kmfOqYedSLTimGzPVZap8yW18S/8ISZFEqmJu62xMAj+1XiInJ37xTM8K+LlMvWVvDX1
/u5tE5H7YJhIWLsfisLRco1FOFfx43WXJdViaElPnfy5TMq9To+dJyq8yyWiWwT7OL6uX1uOZsfu
y1/hvPXjjwPQmHmx/rZnhev/zY92JxsHKmrxjSS3iQKMfxQhar6oJAAsC1Z6+MVKeuA9+jGYUUSI
PfV9wVdrAGrI9o/gXd082FtenGPellsVZbZhijkxGv7sQvLp0hZmmSe4byPoya6fRhkAdAN9Kw6C
Gnofhu0N7nwuvmXaEnS/Q+KB8EC/kR7K0H1vHxPe5w94Tc7Z+UIxFYLdA+AYZ/JJQ5ZjrjoE3JXy
rQLY/4vn5CJPcywtCVGIsVFsdYCAw6/UN/hGxCQGazJzsVyfxM4ULJDjOs9ZpuJN0NzEeEiXlDDF
nZxaIWjzC5dzGgMb5TUMNXaiGcv2nG1uMtmrrm4qXEjE+3jlwTN0T4033x0PKrgscPDDTdZ9PBKY
gY/b4MerZXi3qc5n4fcFt3e++z1O1j0t79vcPpeQWeqSSzWGg7uQ5WSXLZY49yAyYL0++wUtA5uJ
groEHTcgX+HSt3rlar2YaVzenJRkqFeird16LwJ/COgefgfzOcFMJakgarZwn/Lb0WA+z7x9PtDo
dOLBj3rhELfxfPiFQ4YK3zugq7/8rv2ZbMep4Rs8ZwfbG1O1/c6EpnqE8ji4EAEnF4SvhDV1oEDd
DVCu4tHsckLDEvt5YgY2PoM9T5jMI4Z57C7AXffwx/BVSl1zV5HXTbHVQPLKPWJHAYFBiPHHHMq4
zKiEY2zah7/sePqMVyTBBblto6qQEWfs2GE6d+yhcjME3EUMI8gbnMoySnXNKoSpurDtZnR/DM/Y
bMszS/5fWyokeqkezaaXcrCUZjeV21nzMDRET7iKpNzXxfCfkE9J5ijyO0i/JejyBPYHbWUsRAjX
jqe4OOIIuB0m6xcb9kKRu3Hy4oqjFxgsiPXUF0ujZi/FHilnIiw6QN4NfwTmcbNIs5+hxjMsLene
FwybE7LmvreQyCU3H8pCN4RS5LUUHX/iyZl0EQS9QyfBlB8w1TlL06s8pifhMFwvPc/fwQ9ExN0o
3j4kQHvFxf/f0dA4f5foJmfk6be43Mzfi2VbKkKNxOgft7Ql1taQIXqs3Lz0DgWL5m6Gcq0NW3cZ
gs4Grikr39QC0an1ktJ16IfYyMyyKajwhiTo57XzIOQkCMdTXxKk1uKjULnp3dIVA9Y26Sj4k8Gt
o0D9OCyNbIu3ScgTUoK3p98mzn1q7nk+DCaYeNeSX1n90kyiZmSia0+JFH4jBBDsSqrBnqoWNjAq
iE2+i2shpNwRTB/ao/0Opoueit670+IcUZ4wwtBVqtYz+XWtofCY2QBY9KTUp51YcZQc8yk/+BWS
VRJ47r0PfJ1/lPi88X9b0OdWIhbCfyBuJz4zuxaYYbgHQ73NYpgtY4WKtS+1T29tbQpiAAPUe4eP
bdy+V8KUViL2UG4nFoqvJlcWHdZq27nEF0GQs1FADxSRxJRmOSY25qTq2nWognlJ978ywkVZrYlt
VuWR/lNtjZelMEbo11NL/ea7heb9ptuNS1bsywfYmNOQXSs8hOghJOPXLFIUad5Popb9WghiJFtc
bTWAqHm1Fi8hz2qIdSrwJxlLDNN6jpkxp0cTQNte6tuf3/lyCPiTXFB2k06GTQKbp3WDJHoukbzF
ow9Qc6V0ybFZQzpq6BX281nL+Vndpa/j+fxSsEc3dGBMM3I/yhjvUrBGtH6L0GQllCVvZqYbc1rQ
8CxmekPOhU3cx5AXOtwTVbfpTgnAm+7Xuzymtb6n/INtS3o2mD1AasIesQqoDRjMlosAVZ1AMRbr
IvzJBeN8MJYJVvOD0ZfklGKSC2aKU1tNgGjk49E7j4Dbla/9rOy4FkBDDRs2d3Oko8Y3aphmDKyd
RY7V8kJCBONO11OfedFAvpFR91el230t+S2KV0iRImmkH5Q3IkqYv9el1Ev2q59QnfOGEVTC9suG
p9AMHsQ5K9PGK7zNgprcj5h1nGFnTrUXEPmksTlXLdq2iRr9RNncnkWNuSGTFFEfcC4RMp/vssOz
ZQadrMcmPZ0/GW+XDF4SGT9Vh98zdimiqFQwAPWGOhwrIN4X/uoCOxDzK4sptLoP0B54zHeAsRBQ
8BptC6MFm1rOnictNP4KTlgJZoNtbov4JDFzSsojYqc+e9Dip6UAFKRPTP6xEbDuh0sAjPkgbo4n
h2HQcunXLlddbBLuiy98/EpvHaMuUEhXuDX6diFUO5np/m4Zm6xV0eLXbfXC1Uhiu5Ay74ySK95A
43eOMbQfdc9poR69Q7zf8KG7SIQ1LpuonZ7TeCKm9moKTKI1Mjnw1/QZFFv04ZX5wUxNkUSEyDXG
BzIaHQ9VbQNC6caU0bh15/yejdpbTtLxgojjjlKgaEI7YmXSi2i61XXnMafiteV2cdMvp2uyGVpp
qQpZfYOn7YJN3+9CH8VpCnWAoDIYWuNV5GAiRHMvka8z4JZ7WQ9USn5wt0Lz5rb0Hxl1kkBpnSKT
D/+G/9FJgibY/6rX2PYfdRFrxxh0Ujf5ZtWCl++WzgrasRI6L6df9Qji14EtK7uxs+5/4eKRikY4
TYgGtyPjH539pNKYgBha7Jin9ec7zC23GHCwGUtm4YmSMiKhuvoTlA4SHd6gIie6oI6KFx3BOTCs
zky/U1HQ5DZzSad6zPOSJ6ktERV/72LSwpILl3ocMFTucRyoYsZT1cRYr70XudxhK4DmFdXm07Og
O1P87r62C7qF+zzeEMGHsxbKyBJ7Wu2cnra4e5E/WQ1KWSD8OakhecScheXi0ZP5x+TySRYp++ZH
7sQKPVedUPnzYWzEY/bUJYIZZF2UyxOG4W7MsGNcAJT2c5HzAp21x7e+iS/VBdbHQ3qAM3HRmcy1
s+LrLoKG3UOal/aNc6J9jIQfwWLOG7BLVYUYEka4mz07QWv9m62afodEXKtDU7v0F7V6RdXHyyIx
irDw/cvoUV+RDd/DuITZ5Ky9/8GmQ2Ll0nq8adFZDZhd2PyTM0+1ixtEnEqrYvQW6ZSnkBKarTlF
PpdS5Dvdvrlpch+aECLCcvO6lQcRvhMLfqxx5L6FEvwK2pctvSWDJCZmQwFJUEmztVGY9VoZrlUg
iFs3hJp8zNetkaDOsrCTR/Mp8Zq9po6MsFUvQNYBgwybFWXFHq5hglCraNBK2X59MtbefV7Zdfka
4wYbw3R5599fOC5a0uSBH2mub8WvDip9I++VGzgHH1rAUzIh2ibhzyqyH0Qkk3j493BwWoa1pjUO
7+gjE05AR589Zrapf3gXpt9eJCmCV0BlUp2wGd1FyRhpPyaPSO2iDVmm1i4BMrauPB27Ps1eZTXe
ylqBxJtooVpqLiQ8auBfO/5a/e7PB4zIpTROQDiZUF1o4xW77ifLZMYQfD6OdXkDDNfIcQGuiqhZ
mLse8fe7fJXeznRL4Nw+9djyoxaIC9WaVlEiiKe5r1MT9Om49+lPkNrk6ibi6YuDXP2RaAJO8m2Q
tM0s8VTeQ1uVYjzM+K0i5jWeeuU8bn7TML5c6+RYdzrnZ1UKxQFvIjRBCkAAIRVX7Ywedv4l45e2
3pWzRNhWdL8LI9O/fxWlCDBzo2bG/s3vih0TSQ+sKinEesllCen2W2DJ6MGlguh6YrjiT2+4MiV3
huuni2YBLFvzOZpsvC2i5D2N1ojIFB9zikjuhmurhc5JHzi8YMwatqb9S8WAeB1FsmeWXNVe0+YH
kXe2OKL9fuOtRFYz69wgIceqnuS5E9+ORbYwqoIRsOsE2A8DAWWPjDkw7h66nmGMnPNWryWk6QZx
ZOzsv58x0NZOV2CxmX71mQJRX5H/MdCT0xRhxz/V9far80OaHYiJyoh/YBW2jUwPnDeP7joDVij1
Ciaq3STUxKAzRBGg1c6yr94JGNm4o9QSVRfX+DpRTjVdGl0c9TtFa/s0E9U4SYnwyb6ZNipiooNP
kjAfl0i8Rqtr1TF9i5l3RpoCe8ZKpDTpL5bB0134DZKxoWsy3/d3zI69iYUgEiRoISWQd1Wftq5h
KY5KfA6WQmogXacHy++XUI482+3eQn+4cpXIyZJtaqsuJ0L5tHsRiDsRDR6LlUjB91t+I7ix+E/I
R0jRloJBLq79QQ83u95yIAfS10q2fxmEg98h9NsMQ5oGliGW0mgcCFoTJlGiHdrdwnow2rdDB+25
eP0p3FrsEHCjby3ZMM9jts2T8D6ksKesjNWygN2yf9jaYBu8gjGQrH2aSw2ssKI9vdElPN0wRw+P
752mdDcbCljup/mmqcRqSA5EZuCxbcdOy7ohBxjSWv7BlvihTkkBonBwKE73mGJ2FZrkD5Q1Kwer
wWF9oC+YMcC/tfmyZF4ZVt9SYuAEj1a1HKgjklDrwtGohbiQi+z5UyEebCFbO8Z9ZHRA2u3kLcb/
7veJu/o9TspYkcizn8ZJdM8iN2cBZhkqeJVNyHeYkAIjNbgQ+AFMBaltV8t+E/LWiPd9dVbe9Ll8
tqxmRCGdwtxRBM4uhT4RSNu4mAL/wV/0BCqDrhlxBQpUzupbAh3np188iwF8jkhkrG7d+46sENeU
+tu1cpyCifMK7KL7WVrCuBY5kWqCckBqVwaaGjX4G2Nc92JZVR3C8hoDW5OhiUSnCMnFc8wXR3+K
SHPbcBMEh71Nh5aFr9/VpIRKAivoujuK+WsBl9a9h/844RVxSZfQIPBLeix24mTWNQ7oZMIibxeJ
6hiG8XJurGR82n6+Wz6vqNIkqGP3ETqtvrWylkOlBUXt0x+Y3TDLMqXdyCkEENPpCz5mqgP0YBQV
2CjNJh3bPWHwtOM6GKbnKAd8cPYBa31IEWEUBRaP4HYqyQt6/4jK/LdbyTXCMJqZh5p1dOT84OMT
OGB6aWks0F8LOFQ3B9U288ShGT7kFWaYDG4X3+Bb6MGECoyyrBe7e2uXHbv96DaTmRFLZuefLhQl
gChk10BJTnvrdGDnVAsa8pvLaZAYnxuKv1txdiXMmDmHDwj3G2mMvpWeawyHcGP4pxmTyZXr56wK
qfeEMzsscrG9JOf8cgl0reph/6JESfah/v9zytiTdoRQqLAsF8KypTFRo91V/1TTh50GvOgwA+I3
n29roT0v3CKGC7qn3Mcb2MUwwdMJ9LpEvDgIyGvzYCZgXi7KBgXMeGr6UVA5dgXsaW1y9wQSGTZU
uq7ee7l7+cwVh8VdaLxGarFNPb9hO9DkdNk4pGVye82Jq7zCBZhDpgDO4JX5nwpNOCUfaYg+lioQ
S9WUR+izH9Qkcv6sxJwbFWT2P2yPSe8WBBQoymBUZLZDIwUZiPl/woICI+0dIjenaLcmIkGliLQQ
ZjYb7SSi2UX5aSfwPe7ryKAdy0BZrS79mGV7eWdfwuiUwLG7L9evjihd9m0SlJsf84LXst4rv4HE
eIhWqY4Hf6KVQtCG62rmc6SJtRvBTbwuo6BCLrKXLF2LInCNbB7MMHCdrNwl9gvT04Dca89nECZn
7ujx3e7ko0P1/64KXnrQ4Pux9bjwUgEFBDc17ZWxz3n1R+6OzX2hkrdxW++R8t3Nr6JQ4zSLY45c
0dmaLC0tJnqWkHdHb84MxSdD6/iffxuZaG79mkLxLdY6xhxAoHzj6EVPTYXCehLrx80r7spsiglm
Mh7WX+ySPt2tNAAZ2NOXd8Doy86Zs9+TuYiejANZS+2nwvpA3neeK+XKM01Li8bsHZA8qojCWyc5
d0BdGUP/9oFXSmCTL/cYjNs1ZLRxVNyWYxmjeYsb3ItxNYokLh4KA38U3ZfLatJNBNP1F7wU6ZZz
RIInIFi0f8+3sJBcS39/gM6/mxc2Cs/2ohCuGHXd3/307nBgxrYko2gi3v35rxRB4DWfRHHo0JxI
vpLHge7AyrxUB53pPZUhdBvM1oNT+8jh6igEAXLkN162Eb49RbJ6pdjRjtAia26UjIZH4vj/kdrW
i0soX1HFvHZRuhT91/l2wq+xSv8PY02H4JuNSAU9cLZlCkEweB6crNFZlQikzJjeKJ1Ssot4G1MB
zyR241ltGeJgrGMlmKgARAUSfsQlY3AKFIC3ZwOGEvv0HMbZS3Lt6TUIaBk05TtneZtA9tGxgQvN
VmOWcvRIm4XfUHBrt8PP16ZERcNFMv9B/qsVeVuQVx2mm+VwAhxks6k2oC+SlWKr/ZOAqR+H4cpv
iOHrlcvdIEkWN0li9TicMUQl/L1CTPMm88dw+zhQzAiK3pf++SZhgAVla13cQSdGFfmtvtOFx0kV
Ns+AYo2nxdk/LrYwmfkGdsZt/ShkQMHsWmbM/u+dH0O1PsTtnMMcbPctkVVlZH/xgQWFQUl48vaQ
Yz9ZlwpUv6uy38VhINsRSx5ZgpiF735FqwCTOfJICWeVRdD2UsO9bvClfuKr2NtBPAAM5xzQwYaS
h/gmLWcEOzPQO6ghLRToSTlZrjckQzdVFC4kpQgK7BiXOdJPVCuRdQecda4X/v2ERDd2DmIeKfXN
9HiGf/yRio+xw9zIQntj4DPbUXAu3KV9rLH7yaf9ExLvC/Tnbj3Do/qVDRmZmkgB25Rt9dAHdtFu
4c/2lF+nk9dX6xxwQJkEdciK+4VqTTtmmY0RwBizppfhy0GJ/nyasz/MStG/xFMuEJa3kPv54eDE
cckg4rxOTLFarhwF8yGcmvab9eRSDB2wawq+3q4lLLcOWFrNtXz92LUPEvwRJ+Z8jBoGl78laEoV
LhEy/HUFoHMaLn0COKu0cKDXrXbusry4Xbj0UvZRdzd2Zq7qByTMlSDWlsy6hrzZa+nKoEnqg4mM
IOXmzrhcUi2+WIYyLNWs7gTKFxnP5bwSCiGV32J6d8LyiAvAQ3OR8ejNw1Uwj0YKbwNn9XAVSo/k
iJBPk+Xc0Y6oDe+cgd7MtXFQIFQzD0DVhmqgYzWno441vsOX4s7PGsy3/kljPbGQANeRLR4dX5Ou
oi+deIgBaeXNATppMbtgrt/YlU8OLF/hRPk/OnNC+LeR1FLcc85ptLE5b+EbO5ItSa3u5kRc9+Cq
vV+PpTnO1BYBgA19ss7oR0lAp1qbSTpgiixK++OVbSf3VRviUFfr8awiyvmln1oY6KuLvMVj3pn/
NgmIPduGNSuvNrFk3s283o3Cj7f7F8TSZC99J3gIblcnh7euwb6P5qqNXoz6ohpU5F9tbq0Vn3Pk
QUuvp69jqDDcSZyOk6ef/ncBPLfPQo6jFNOB3O3+3vFqRY8uCgCgba2ua/7aXOiDFpnqqn22zSIG
9QwfAhMWR32If8XDtoPyex9VsL3lTuiSB45tH3vomi8ucN90R3rymnDcYXF8qOy4Zyj5GpJF3Jg6
p/5a0YIbDGq2phAnb3HKQfRjhNF1z9hXSOHa5IQV86p24ume8/ctt4K2gdfcuReFGb++kHrPMBNv
k6b7USEDKN5uJlSWZbiBgryNHnkYLP4nmtToyUPLBeeUL4pfp60ccmsNNM2F+b7TrCnd+Vbq5GMv
J7E02FZLROSdN79bFPGJqluGWsmzBmSx6RHEuPdLpqjj94/bYmtgE7ERId2GyLHQ+RopUxEUPUSL
/bVRFAKTraKw8H9dLU6JcbwIcMgrFzkonS4WkrgQrRaqRh6L68IViJ2tNXI4ZPZxJtYVjpI+XulN
2sV63uQhXH9mHKm/6niSUmmUbwMatB/z+CdnCCfDolqFzx3f680kbee37QY/nqTfoyDZgHz2r6kd
4XuSxYgPg3gE6FbYsiEMkpAHA60pS2pvkrZv5i1jeTz352GIvSjaBajwVKNWh8zveBHREunI07qU
lx7m+SbfWY8yFgpkcbQXv8qiCGbb+WcxM7FH3X8Hce+IH4vZPjZVucqiSQ3AF57OMKK3eR/tP2d4
h39MGheBHqrdDPZOyhXb6aaUFvbGXRHEQvEA2NO9UxzC4pV30Ay9qeKG89tHiPT8/M7JArPvvSo7
vnWdC3DUM423mcI7bhWnnGpqzauRPETl7gCydk2hpDl7Kd8qhUP/wq9fJPy5Aq5lCBQH5xqqSlov
asPrNdfb57wZesgCvscGJzf8HotjbQxZVwDPgh0klg+kCmXwmvmzrU61TTBNNy7SeoSBwVLKAgpp
J5ziVdfGO4Lhl9sudAlJXli98LmRHF2MvYw4cQC9I6bOAB3Mhwk5laIhoty3WpSXunRyzFJWnpDa
09285IbFCtlv0Xm2OGFR/XExw0gIOa84dRyAGjK+ACN7Rz9YkkZj7BBiTQz+uU3kJRVA0KgeBGLz
K8J/E1mklacYjrW+lYirRQQJppTPl/b1qO9v8T3I1BTLUJVM1MZKUHYTM9coGE/h5KHTYG1vhZF2
ye0rAGqv5L0qGOl7FddCETu1EU80ZwGYLBz6xe8v2zf12sKQgVlW0qnRzr2ik+33720dnB2/qF+I
OyFF6MC12oIl8kEAZX/JAtoHixbRGIJpDsDhr6ym7ANNq2la8nPQ8AKifmLEJXjEeteYd3zRnvs9
n049Pg/GFsoGllLM0HBLXs+hNr61lsUHth2muhlfn0I85DzeL5YsNYN5N5ACRGQ/qyRz86zI1q5t
x6GlKnz3k8t/ZbhAkQiBocQpa0oUI+TEj+HUDnuF0zEmJyQY+guAjXf2M2UT5LDy+q5iHrxQfdSb
kaXPpiqD/ZFA9ToEqTrmwwQFeTZFRMcgqQetG3Mi/Fo7QvWw4y/WxejeTWTIliz7tDN7Rf8RecVz
sPNdW/F4XWaw/r7PLELsMyuPN4sm+RSnybVXVEClzfI8xLGbpNxfLDYmhz0+xt4OHb/I11e7qNGr
TwUXwvMWzGaSizKX2kPmwoBRUn57Oi9lijGjo72k0L6yox63ADRbSC35kSMIqGX805OtMO+pk8mV
0Xa9cSAhfEjG7HijxeqrRNR5+WVDaQKnigmGI7zKyH4C5hrG7Jfi4GNFRDQ1jgUP27AiOBn5pKLy
FNZURoELWGR/CiehLTDYWHyT75XwWlDrCJmAX7C1E0JucewwISm1u88t6Hl/2NrRGXlk6zsaLmqK
k+2q5KS8Uk1T08Ckrt0qbiIYemp5ZBfNFCYAgnb3Dv9UBpT2U9mbvbXADD9lBhbLxpPGa1eQOmyC
/lvW/m4p+DlGFiuGvwHe1XuW/RYcUvf7bRyuJiTRjTVW/sqncaayftVdypmyVHIc6b3DK20tnku9
8u/U/LJUNxSyyicOAWv/yjKheILAB8Y+FOEisysJeoYLTxANFKqx2zh99OuP15cARk/lz+4l4+l2
yS3/3WPfVaxueurHOm+Rg96Av9tVof5g0fUSc00xxEWEQey4Iycnjtz644dUq8JskAZjY+zANXJd
8lxs7Kue3VLSFM60/nUBmYgBM8RNwi5Ok3u/0T3xXu6DDjaeQoQ2W/WjIKhqb7XiawoSkSuGxSje
5e7FA2Chx9jgUnrhOUXsBC6wdArgUdVxZxsFQBLjy0rydOwS1IPMfXcS6kG9kk8FTHh2eu7sF+2G
aXWW0FBREqW6g136qoV/pUU+BvWH0xayfI7WPxARB+GdsOhuBl+WX9kOiYu0Z6icGPRUba48Aso6
YFnqNgc8fkIKnwueVeiIdQNI1T+85laOTrRtNbqiPvUxHIWwCBowe7BCiiftfVRkImTFIr0frl79
QXjLiJ0cOzzoGNUSK58bl15e6Hhb79sDBE8ZVzMVr2xBDL+6eAoalvruJIv0KW1QVqnLf9dcbQyk
PuEDHtFqEKF73mTmV1gPf4PM0tKdkg8uK9RO6K81jUoYb43lArXDM8Em7X5GJdvYrotlUeqXBN0I
WvnrJqIGZmw5rHHNqv6FO4751w6zpp/rwXUKuKn9fCwCieHPrp/oS3mCnAGb1VttyKWbE4bNOQVs
CasqI+m1CW9QD/W0gKZRM7vykb6bk20N6erETC6jlX9TPBWii1p8UteSlf19IwvX6b9Vq2zAPM48
jborEWy8p/aIMjJZUgRbr6FJ2OCTFWFIWa7p6Qb4jXRZTyjWWpKn8intuqNe7qZZW2DUzYxGeaTb
ma6qPTlONmH7BJ4t1e5Pop0T4JM8pjum4xzc6KVhs0MHSSNrdI+YodwYp2cg/stz1j6174I/22yC
2n1PvzSjAHakFRtwjAtIMolLNy7BJYW/Vlp8Nb7v/bqBUq1E2YmwWYaYxzQad0gxuI1+hSqLfQeQ
oDAKCL7cvnC24XULOHxCk6osLBkRaShKYPR11Htx6qV0zQHf7LdhVE66eZ+B0YgNHzD6lXkuYSQU
ENqtXJ3ZSGrkFd1eaPvpVEPrtqyV/AqYMEKztUYSjEMlyURE0TUG1yDvSxjkQXHjaP6ubASw5V9X
/vgbU0lE6DM47FnghpLmIM9ijAtqcgrRIIfvXp/U5c5j6dFLthKoMVudgVVBO1ULLiXGYebVuC0Y
nQ4tJHbLDZpIMge2dUMWMWSAspHPLaByQydG2Q006zBeOqWgMFlsUexqKDvX2q2ntmMhThoaKB3l
6r0BV0OBe3FPfptjwmWMA5hF091M6fhspQjIcMtbcJ+iYCs5xsIp9AKo78Al4BcX57yplhWvyn41
rTHk2Yj3L0mWlLAKO5hkKrttIMkfQ+qMnIaCG3BT7jS8hn8BMgiW0NVfgIJf6DsL91scFAiwZlE+
yrTCmzdyb3YjePjWJN5wnv985yrX0yY3ZRqkIhdobT8J39RNnWUMT/b6Z7NwX+E671zkS3GQlT44
855X2bnneKMyA1hBuAuUO91qvUQuq2hVnvuItgDf44uktcRo3Fr6+M7POiHs5d86zvRBVtQL0yTl
BM0kXNeV43uM3SMqPMAvgiWCK+nnjw1ao75y7ZpCS2uqTiY86HvOAMJ3IFqThp4u3xufYj4Htrlt
Qd6rM+xPyy6zg3orlgU8lGefPyjSKDFJYws1Z73zajb7YN2YS/mjgm5/voNctYi1K7qMwEJgaW6C
2pow/lyBy/sfXef0CoNszkrld17B9lA0LCXw9rXWvEO545DSlx0J80GpfCE7fPSkcOt6BpXJNzuR
9P0k9i/CFqFzONAJcQyppsO3TZ3KkhAEzS3zw8Tiw2ripueaAl8+9nAVOB20Ju5y3SgBZMnxtffV
BqzW4MyDku1fZIfGSvoRpusVSTxwZQJmKNrm4+6+ZtIiKmJhqxoCqm9jq9Yxp2ATeB2286fylJv2
B30HkfT0dTlSDeeg+zuUPEQQigStpLyrIPD1ErjJjM1Q2vGZc20J/MNGf5PGzinkxPS9cx+gj085
mPywVdPA13TCR02VddrajVB9fPx2G6NKYXgBJpvBFqCzqdh64Y9MkbUN1TTpYAPhb49+NfVAKpql
U8cpLzdQO3r3ekK5LN0pf5dsdvUDsigP8L56z2QLd3+FqbB4kUT74LLwCQLCXmfCLp5xPVuCXNAC
yZU68N4awiiSr5h0fhg5zIqx9L1TbuHV9R4a4zYHPMpA1Pf10j2F5qlC99E9W2+iLd95WHx5zg1+
GMv4bBpEg5k+QP4QK3mu4z018hs5plOsBqvsE0XT661jdOLllYKIvqD7YqTopkqRmufRjVcE38FI
V+jgOrs2f5uPI6tU/ULL8hjoOnBlJuBeOQjWOOlOlfgTYin0T6fTRs35c63rpSSbRk/vSabtfQ3k
41CBFxqJK98ZCH0kfirso3mMdWcjWbNJUilXogyrsH8prEuWgU2qlcRxnBRf4caAHtuCPkJsqaAh
u9ISi195hrr8xSeO+lACK5eCfktRLQUwWBGg4RzlkmOgUu7CrFeB9UO8AF6UkEYkjLzH1oUAoYQv
P28dpGGhQCbRJSQlp+m2mIvJ9XJmI0myAFp79axLbh5UpxUz3ejaWLxdMvfExUQTWRYp791JrkwT
pfa1gPJhslsp664FG15+cQS+CKpkEZJxcqoTP/LWhxqxQ3vR/ayJybTwUMOrDjm2eSYZQtrNMWw+
lKGTE8JSRjIBHsIiIq3fMhdpuez5mheSQgXjwyOU+IfGeHhvfsngrGg6TH5y+5uo+4UAFi+d0Ttr
P7xJoIartIjsJG3WDGuJhW972/CSiVo6tb1uP4TOVT7AwHkFPTfmxSGGDRkRJst0J/6WA9oGjvX3
YPc4OwfYVcT6Je54n7sD6weTYEgSDM3ybXYPHHRyreq2lvnuTC5k5ZYoigNunH0YEcxiY5Qm2sL8
MXnZlr3EnErebEgiAEeOVbX6FTLeRPyBJiTZT1i3sIUhP2bSA8Z6arhK++JigxOvXNYH/HDQgM33
8h/gVxj9j3ju0CsS5VsMofQK6sNOeXXNlOjMU+SxXpzFBqaYsbTXe/xo+VMkQZXk3IPxMFe/VHdq
Gwm9xYsbpxgBbFkk6qLVwh49t62MPiDGPFuirMQ3chMjMfQs2R/CSRBTPBSP/oNdiHBJOCVWoMiH
rweQM8xQwzf/rZa6+DXFzCV//8CPTpOXOcO6C7b6CbHt/7+Hr6YdHA2MGfWon+vyaWTjVyUNjNYf
F0pfRLObAo1rZX4imRFiJj7bx+mUaD/7Lx4fR/kX4D2W9Uqh+WcLOuULEBGdjYBP347dbaoAAyPl
iuYePGqZYK/H+0CFJG9+/KZVAUPAR6deavPykfJzeXnaTJjrNcefz0ceqqycvBmEjjiZ0/dgya1t
aZmpt2FVOi+Up+AuSd1CUAVXL4CTBQYZSWQrniVD5XJV5ddi2NEcToOaI7AnDAbKlvmal2lUXDbT
cY1SmNtTNcPLy1WQaiw8gKUIvoxv2kgbNv0tovYlbSMBf2/avBtL3hl+T0t9ORiK8PNWARLS9h4i
4M+N7+N2YMMUZ0YBfSrx/9s+sjQD00NFm/muNwJpO5Q4H38VEm++nbWneKg8qWQpkXk+M458+fTr
4cW5cKgYB+fICWK1+M0HYcDR0GtvVhnysew4PfbjPcLb1PeAyCL8bgu57J78l0hkVMqmHZw9hzP0
XWOxZSrKsP5+28BcPAJWlzkRU/liAzbYK+HmJ6SRkKyczd+bklepC/qaOgtPL51K71n1YKfBUzgU
V/qzHFdOmO3pfDM+IvWhvSrpJN+CH1QPI0ZXDknPES+ial1QwRIuh3c4K1OubqzTV0Onx+GCjjRm
PYnhBcA367l582Y0wB1PBUhuXIBz3HGbio/rO/a/i1f70zykJGLIjM7WFuwqFkFqtxu8y+LWbHyL
haiQ9XxJ7HDczT/7wryrIR7jvW1q90tdq7HI55vr/ZhQFbA6MRncpag1ScXib3EGg6h9SCeu4oCi
5UZ0JIs42kZLKS/nnO//WmkRglnxd5P6WUAg/d7l1gLKwv5twf7ZoqN80htUY/eIXFOxBajbzyGo
iWEmg55QmtZb96xaOtquQKG/ASy449nqrpV6U2a0r+FAD0/5Qw0WaiC8ZyuFmPVRez0HG0+Gec0g
zQlYATLIbT2jlbHhwLIlb6XFuJ3daak02kCJ62iLnIG6mLUOvnHJOK3BhwUf8HaN2Cu0YGgYMc3j
wcCZ2oOnqdFvrCTeIwrJQaBpFVAduZ85cxChe1FpcwFH0hbtryCoBArST0lkRNGLpu6+/OhKPa3o
4r5W24bBIfdf84ALvyKYmJ9q7tGsfAtV9THgJfbe59ACZxh/rYRrq0PrfFBVa6iIuZL8sYcXFuAe
RII0z7pA30jb5YvOHxwH8GeKHf6DbNJJ3f8WO9NYVDd8FrXAPAw5hqrrq8PP60cByqkR5D2bjEkl
w8qJ4p1wIgwRxq5jguGT/TuL564iX6EUrKastYjxoJe6kIWCzrkg3lsbTNFXGpCWOqB0XEV35+Q9
mOOd0YYPf82czxHX0jcAN2yDaFOug9O+tysdnDj9HN8aE4XS3pujeHpgTUg3WzT2w83BZ47GRkCn
F4hbxJ8P/a64/Yw9zOzX0mjDVe4e6v2bcBoMSE0zaUrzY7eUj4/bm8CfcWcjaIsQaEh7oLFEUqxx
yCfk6/h/xhyHbF4V9gHg4hYWoNmk3xPBNDR6hkHfk0Mdo8sTUPuhOyyK4OUKixbUFvcSJaLlhom8
epkihfd2UA+O180TWGWyDfGdEGMJ+vy9wl4bubjiGw0UJN+d72iusOJfpApOL5TrSFwnvLLc66ln
eiIWk4S7NMJadsdoLl8m81i8meJYDFxA72rFpoOJX78LL7v5nj1IgnC3VFepKyBzfnOUe9+h64w2
GvcqKaICXDTRGbpL7avBrwZxCr25RTTechf5TNo84f7o9wETa0ZFZ7JapkAACRAYMbysUzn3YPHp
ABErNkkVFR24EZ9eQ9GD0XLz7/ygxgvGBbSTCaSfQ0XDhj9sYJ/fnqjE8EqmL0ZIfQa9iWDjxOgd
qK0bxPTbaeDcKPp+sHpx+FmnRNyKo5zyQOzQiOLygQEk6Hu+pBJGvnRXp2oJH9VJk1aV+ZjF+5H5
Hdxozm8r2j6e+tjbU9nBbYs+LJz3x1OfXwYUJlKg/sItwLcbn+YlDweCutxF76Cb92uLwNCuIXA2
1TREkAk/+kElvxScLCmr1A4ZXhbJdXIG4iqazZ7eVn+5b+co1uTTIfRji++1VzD3fECgeVBueQ+a
4L9qNTUJ5l9IfLqxi5tymaWQ9UW14Qggtf0oSU4AJ1yUCIN9/oCaqqdyk5DuoPflBP8FpGT8CBHV
X9XhWl6D7Sv9yhZO6sAiqBOMZWea3gTf3aSyMIZDZpTIKj24QzqJK0801c7d1qZtFXHCl7TxkXCi
WSpDLXkjBiXvP8mi+5FEf+mcfkgZfo+PiN3u2glGpEWoqalSi7NZ3ThPbUPhu8mfrMX79ZE9dlk4
S6VDwLJ0rat/5SHMcJUSME6OP944iFey6cw1eoSBfuPHEGS1/PZ3N7cYOL2J3eMD2ox8hC0G6hnj
u1ZZ2X5cREcUSJt3/nOfZ27eQadoIVGimIY9ZLBtZPiF7K7CuZb/JoBgE1fWCu6e9krO/xNZWR4Z
tNLgAaozPoripw/iJ/C+w8Tsx53+SuTheceZoFV6vPr750PPKcExOpBJSPZB9tI7MYd6HVTrH+Yd
I6KYHkHerk9MsgI03RvTw35THI1VIXBABrbZWe0P1rBHxRS7i+DwfGhG3ct/bHr7IF/4tRixMuWq
HkUj5U7PpzOsVoGseE29c2Fz+S9Yv0bSGsiKNPMwIcwPmTl/q5LPoIZxfDDmrzBp82KwMSmfapkq
Bw8gRMugavjn2ADAPr8PZHTbkdrNSgDT3t5yPjFMkwQsKNMApNUyeGnUEXGUUgKUAJB6pUGVoJrR
phsuKV6EoVSiRGYz+9J4ptdLytV0s2wlwTvv/SahPYjESk7cgQvuVjq4mzi+74egOIr4RtJtoEPC
uh/a+AQrdxf9pNxd3KxC9UXUFP6GshwG1fcBBHJhKiz/uV7B1JJQiRNKNOH7becH7CNtjfoGVMkX
hisO4nSqRBACHvWFRbVU+3fiJSnRhaiUlCfqM5Vpb2CXrdr55SDPKE1nBhUvD/NO07BQPnQRfogK
I+4K0hnjS830H0VjJFVAWI2uH9lVakBXwO7vvJi6jZRcc4Mq7nF+eUP7W+EB/UYObP+AATLPAwxD
v6iHTT9XKsvwFWJotWxgO+EAWcZ+ynH4M73fsOMlBT5DpyWo18xaH/d2mvn2O/BtbqTmQFpRt6lv
DkOMndPlfsmDTQWw1Szp76jwVTsrY5RHlN5aM4urwe+hV5jCqMSeUi74RSIJ4ca6Nf8xjwDa+Nd4
Bazxk58B63tjX1rt6lml/vtriiN8Tw2ncYll6W/zYBci9meVCIEKn1iLNnjsYNqY8L+u7YZVvIU6
PugZ6qOVq0TJRp/RfFQymPLL8ezH+DOz1pPf6Hfmpua/z13jKdMLbHBnpdLUPCcEqvTCXKeTTgD7
qhYTP2/X4mU9DoALHmab4F4LjKVWVV8f/3r7Ylwazw0weeb1SyFJ+QyAyjdfaymOwhrylijPtNsh
FhKboIjd/vULUbChfQleTgryhPdFjKkCB71O9tc9KX9psAgbyi9RDUf6Mdf5uh5G6Df+Dubd++3v
N7UntT3hrMTP6kBbFxB9/v+t3HRMd1F/Glzfampod6BJkQcQqrgOdBd8PCPck9pTkkacJT+fbQv0
W+iPsodQ4juiuwSncx4AGc8nPsgv/+pX5RMWzqd4suzxT+cFHO7vAQam49WQUnlQ2SF6rpeNY4wr
l98k+VkAeuPkVf5Bfyq692vXOYmMl65cpKoFmbG/+BXNktyHTkbzIUtkYh9iPCjseO+L/gkDELKz
2m59x87uU116+w9BExl2DpZaAPWwCdQZpM3Z+X4gVO4JlOhdpiH9nAYnawe5vSnJzdBrs7Ftrisb
gXiOjClLKu+NF4JEjdJRaL8DAGf6X8+9JMHOZzrWKUbTggH87aYe0jLzuvk70AMCMTCEci44HiPu
4Mwv0+aDRD7C/2vAkDBJHNgm2kOKeOzlscdKyaDRuAcEUdTkTppgqKBlUPw+jIKON9+dJ8dGdO66
2ZHyxglYVg6+HbOgBcaQrP8+K4c/ha4mqeydaqPktZdLOt1Vyjhbc55V8oUPCtrCqxopBu98a1Mw
6sVbNE9BhDrJ8g+Aw5drX6lOBWwQEa6XO7HHLjayy9UvXLa1Pia8kG6hg4YHpgi4Gcc9UTPhbqW5
sq4+XaDtd2Twl1u+2v83Qe/XXBMZ7oTcvq4Mnhl43kb91mkypGZiZqHcrdNHd9msBhL4gpH2rOZm
ApwSHq81fACWz3/p+E3mXn51TMgOH5aAB8WB454yvPxalD7hY1+iF/pzAF33xsF78enNQkagX3k0
I+234297amwit51fE2tC17fASf0gklEPkhO1yuSJP0lcWTsSNFef92qPDcRxkoBc3XE/xWXdGedx
LcjxLsJAz+0Sq1GTvWPOERAXDD1Ky421RIEhtZBbLFXtmH8hrhjjLYIdMVz7flqkulL9ig+wLkAc
gE5lv61vrZM0zyf+spgggJfXk2opNDiBU59m+oQ9ulgV4f+40ngBqFGwrQH+XUehedW+lJE6eS//
WeFtAqfzjNHZpwTpVeEi+Wx57znCNrMkLm/+FjCQxN+ISyfH3LYW8lVvpjcIS3bjJdzXSBNcOrwd
ajc6UhOsqWuWNo8IMecIRbgBQtaXV4lzBmdC1CL5WBlS3g5fkZbTBY5eiHu/AYMdeO7Xy9U0DkAY
B4t33o/jA/aOws/nkhe0TW+s8Fojy2oWO7w+0hecot/o56Eulqsm4aK/sSoyi4i4OjkpKOBz7sM7
HSun/aJPTTpj6AsUusLTFI2vEgRDPzQQYnvQpLSO2tFzs5pyKV/q5++ud/W3oSyGQm+tUwe3HBLl
W8qTL5Mu8X10BTJ4cxpE4zfL6T7hi5y2zfHsWs3cxgIJPY03B7rWDionxKRzU4iwEPols0EQZdBm
SnxF6Ne8H66aLiqHwl44sQJPWLo1BIdkkFF7/d0aTN3N1u2PrU2R8osyAnT1zRQZ/qLYLju8wOU9
lp3CJovVmFoiP1Zz5JtjkwYVptO8JTTMEq00h6C7wqHG+mF83GA24e0q/Hb8cnt1Y1ABAPfOH69S
c8PkEw5r1tEWhlKyAIiiB5CS9bBUUlMR/rX6602H6kExdF8fYUCHNinKaIW/9Ye1HjjlB6+Hwnmm
n6FY+nxBBfL5qBWFUHN5VaHjFgwgWidmImlvE3QhLVEQyvSNLYfWPG4+zz8igwOO4/C479mJqLx8
ihYqA8yw0lVTQx6fYdx4D1A9BPGvA96g1dTtChgl/46z2+rVrCj+mdm7fbjZbhJ3wyRJy3pB7ikz
FgM6Z9ue3Uti/0puLAkXywYhUyocmPF1SWkaKEFd5YMGz6tPGyKV2mG9XO+gGSlTSFbBBeSOpcDU
5u/+533CtWnm368bBr7NbGXdkq+JbkKlIm8R97CeDeONwusHHF8g0e7S1bm0iMmJxQ6jOCosaBZ1
/b74Ve0fgJqIa8SeWkhtI7tST/ttN4st0TmHE7akcWVXCK/i26sXMZa2XjZhvWlMr6Cp0UAqF/Lm
r+zbazh/eMz/p56w8LLDYcvEqwIvv888LecK12Pp6UXLhiXDzdXg78E0CGa0NGdqnhTEI3aXfvjo
nN+9BmJ8+xEzWOL8PU3nj5fxvqgH/UaLHKzRtrWLa+ps3HApRQlyBaO2tdIuIEXuHbZb6R6JtS47
3/tiYcphCjodynl0fAn3OeuC/b7T/xCZ0loK35daN6ycOveJcFTMIKmbCCGzz3vCOdtC934zF403
5N5++ny5zakApnrP0nsT7Q+6hst7o2HiZe6xdTfLEvZtnuTfoehjIRiGa+61X9Hbk5m6VD1pTxJ2
HLnT7O7NWAG2aPlcKErgN1HM0E1KeeXSIDAHAOfRUb0faIdUNdUEjNkK0VXUZc5ynJBS+sVZIsIV
4nvSrRZkC3Vl5QV19XaDN6z00F9hCsO9f5jQd5iHqloTWV2NGzbx3f3c1DxIe71qT1lb1SiKCG5e
tUdM3zlvM7pVPqCspOTJyg3l4TD33o4GN2sIXcQs3XBzqDdn3JCYjmf+IvFO8JC2NrtyTyETxG7+
pzUIWcihEI0D9chxQfv1oeVjiUMPcNM69lW7iL6GHz2W2dHXYSMCrUONGEV81R8X/KGv0EAb6PTh
bCuFf3euSWAjwy+tvXtd9539WpRxhqa1yzifQcBcgMFR/JXjYtCWpMsf7ya1nap8oOGy2OP8owt1
RVt5XdhqFn5XB4H5pIwUcVMuzi7gpQaN8JPWJXvaCd/ZQBYr7PoiiOVWkfqrYyk7sIOizFA0S3gP
sHYp6dCkj7PO92PSLAI5dU57oJOuQmN38HsJgjP5hHc7AWUNO+UHGI1w/WjeAHVnhUK296w9UYtK
JtsZicjM2h1wS3NL5/+MZGPPt4YoQqZCy3KGSy5y0bs45200D1N89KNKXU+BOlQkFIDfjV9cxHlg
zEs7bXlAyL44ZErpJnjGTxjJ9SnGODEgCO7bwhktq2r2Kyx/SdVEEV4xqY545dJPZ8dtdFMdh4Sq
+AQREN1HcQ1HFa74mCsMJcN5ugOxyN8Wc9Ly9uM67BpxbePVZ2V6RhusUF6t9mEx1yJjECEVKBRP
gSgLCtBXtvm1sNRikE5SFP96c3tkzyoMF5436mqthQ/1A1EvAgFOM5Y+uQ8fU9Zf+DGO7ysbdKot
28pq8Anz0xh++yACe5Ja1l22NXbfWvHHGKG1Jh1VZExMtAPb80BxA9tSJhpxbn+zIybR6X8HS4YZ
D3hNBAqV+ZC1lWgz2HOfl0MFcjPRvP+mxIE4LWXNTsUlsqrKmqhuL8rbc7VkXpzHiJYThS5hGjim
EIrdYNFjFlqcs4v4F9Bqaa8MZTrKP94gx6dE9aZZF1NVN/3hJZDweIUap0hEPAEKhXYv8MBah3fP
o+2rcJ421bHzRmrJ4E+f5TVKHf4Qlc6E8UIOXjlrCnjJpiT/E0M717C5PUbmLF0hI9AG5EsV9tf8
QKRYI2ilHPJFoaOOTaXRRNcxlXL3ws6zkXSOwrwIQ4haqYFfF57dy5LNVi6TGr5yncTrVGvjKRtS
rlwGK7oOCo5PkZv4gwCKmieluCXHsG1c+mMQkhxK5IS4iumObvqd9xFyS88OhKLKX3MEHcBKyIAk
dOlXsFdP63i4B9yKxy49Gk/DKHyJLwisi9U8sNy7cLSdLgOP/bRcnsDHWQONmonhKwaScRCa3pBD
YpfUWe7J5a42OQieBsRrn8mBeq6zHRzhmsxZSWyDySdOFUvgHjZZYSIA50xskFyhIyYsdas0ohSr
qASyDAZDBRKC5uFiWcwEnT1GoT5bXKDfpuTBPRwctI3keOGfPDD9zVqUUzO6fjM9zIpGtzFfU4hc
xfoPQUql/dBNgxSr52SrjLW6VGnkA5It7O5CPAahVc1ySc+29znMR5MpQjRWhu55iDreqhavL9C7
CnS/14F/5T93pmOyqY2l0hbOJMQk9dc9teWRZbu6J+iqYDdwyIo/IJbmpAo+RsX+m0lF0n/aRS7H
EtXqwG2D6BJfE0JEJIBGsElkH4H8SNjzPQePW7jFxjN/VX3VyUUymC2PdNKmI41R/g1lyYyS+Uoj
RjDnb781280qn++VFe8CUU/rbGkWWUksXdJ5oXV14r7YIfFIl5w4gxyquscbfodSv4OAU7r2LwKv
0e/xVdaGIPbyxZBkq/VwBYvBLo7HmKtu3TPrmM4BQPWO2YNWykZSCZJ5DK1qZLLgQokFsKsAR3W3
XqNjBBFRo9Y54cFWebVzItfA8lf2G2IC3iibHTqe/Pa0Q5sBypGl8Le0UezDDhtFZuwqYXPWV/u6
bAwNVSkXvm+3HuUt64V6CW34ZZFtEduMd5jsMApJeC4JOCrDkTtRFaQj9XyzygBLJ2KRXQDsW1ie
TMlpW0ove+vVaCFdmjn32FODN3sUTAkWiR28ryItoRIFprSryhU+lccJboat1o1oxz3e7wMot8cv
Xm6V+TidjkH9R25oR6Zf2KtIrD+vKgg1+kpPlebiUsFlTTdRtoYzXSN8vJozpDk9aFy2b7Vqk/23
je8k/BlsBEJ8AJItASY518Iv1k4+8iw5B1W0kGdlbiYZUpzD6UlTBpXkw63KDYSyj0sdoWpn0mC5
/LI7PPYbYyfHl9ErwcQqEdyrxyRMJwFwmT9KUO611NnN29zevVh9QTX55ABMBl9Lekf6Srm8+iNX
/Rd2tozUsTlMK6fyLtmrT7IqvnpbqRgGCWig3fXwNSrfjH8TzWlNT3UkVwurfid1mpo31xfZcssB
KT5+hY/N+pXtkmW3F/y2A2CRET1HHPnytgJ4tGyOdCUJBnpRUI2aYHPtN8kbgyYxbyafNXBtOP93
wPMv0GgOZrsT91fV39Jih7HodyDdlCWPIi9YMpx0Da1X3q3q4Z1LKXE+JFNL4QrBexWXkiSmzs/t
L20AqZjhLKEOvvwgJuaaYZYosXdU+rpMV3kYTC2SJbItHDfXQjX96OkasY64YhF9Mi+Fm8cglZmD
k7BosneCgALWdTaKOu8+LQWzuOiZbkqiIywNAvx++ClPg+uOPMkyGdFaI6P3IcBxG79/KPJj8sRP
7l+NB1hoOvUvos5hiD6vLDCHQSAnMfccA4MI3Qiy+YHWukSM/cWfiLNn2wW8B43zd3Hw0wwBdXeA
zF3/wMIMQkXzsf4NbMVbet0lTu6SBsU9Ue2Z1MagfvpGUGtFfQZ+8iZtMWjXL2FKQ60O/oaaRp03
9vePn1HHegM7JLMisJ4o/Vlhm6Fo3bHkX+rgp6RYxhZuEXRn4ijNI7T4yjHPoB7fDbJEtAUw/jAM
0zW+ET0F0ahO3LJLlsAFpct8hc0I1afl9iWYCUiLi44Z8cZJUXv8aXkmZW2uWSIcNfbsgFT+agXA
ODfdMn6vGDhghBdsV/upUzehnWyEBc3+uL/FUxy7aLwHPuaA81QWSeRozoEq20mopsBWWlKrIN15
7T0ntRrw9Fo1/oP1AP0H/HHy9uTmH55Nm6Efn/tjLHM030ihDvfL8xi7SVvLTeZffQUb4YSg1KP/
tDKD7ctIN5ucNM5mOUaNNpVpO8A0hjPciZl51+ZPu91JTL/uPYhikGJ7S6jR+TiJPZp9j+3fPFd5
04ujnPab7m2Z0zk97a6ZdJjbaX9G2MOqGqKlGj6bFuXQRMms/+jUZdlH3opoQ0DN1Mctz8cRdTbW
E2yl4JsxvebEayg462h3/6FyRGjf6PtXaQ3PKPJdYoo3702VPGmPMTiuujg6QwhnImSFKm4dapJM
uEMsp51rsvHQGd1dM3NOYWymFff9yZwNYkloEKquCLwqdExOqChzC/hJTx5akPtEIcExLmxx0+ZR
LuKqCHzr+tll9ydeCg+ph0UZQDK2UOG/0P+XfL/SOho7c/j8bB3C9ScdvH/GVPyXpKvbRnPzu+Hg
tWC9TfuEcV9uVSvI8ZY3ZxUFPfsy2pR9t6BO8pae6FHICleWsMLKTIFLSJ0UmOoaofmrhpQcs/Zt
1ULyweEs/vEGVogR6nf6D6zXt+r6Z1guYOyktaUftdF/4tczgnQ7bR7mfiPJHBbTtJVdslg21IEo
D/s0kI5rymLXPT7r2IhfQikDmnvyeWwtDHL5LDT/aGHvQr7B6vsCGj2rsE9tIzKXDJg2YmOGYy0t
NtVDmq4+pdSCvjD2GOME6Gb0O7c//IbLJYmyycVt/oib+9yNhB22IBuaDrvyvbqstdA/GoIZWJs5
6yT2YDlf6MvxdAky8PyCcaLoqU20IoFqmhHEc5XnsXOGHQlQS73OxiZyBlQHf2MhTzJJH4v2CIhN
KgnvaooVh1WJsL/RudmuVb3UITKYDOG5YlBabDau1ekpg2IbrhzXZWPUMmJaRt+AZWTkf+cnpXCC
CwJpFPEKkD75W/BNg5NE1GJy/YFG8+0i0wDwXKTMii49bI65PdF1nwGZHTcKihjF5lSLOOak593u
NMAn1QHSA9/65pMHzpLiubCA+KWrwAmZdFNpFWNmxgmIifd7/ZnGMFX1H2YBnwovs/WjlWTEYMlc
5Ibi6DU6mYvBsSxOCwqarrnottrH+XrYFAbsT7vv7t8NSEOYZ+hq8vqmVn5UcZat4qOOSg9+EzzG
eMB6jSvLyNlUZyNll9a/MWfHg3YRWfG76HMxcdOdhaNbZn1ffMC2KamQN3N0v4Vq3YMMS8grD4Gj
tMyDKqALNLdigQq5dawkXqO6gyynK6eX3apxwyydPIymPNWt7SgWIQTi2dhVu6o3AED/jZro1J4J
PBDgAMw0DHWNclB5fuTrQLArJa0p7DwZdcm4i2nfpa/kE0D9xSciSjY77jdGkN5IzgbKgF49Cg5x
QbHlw+JX9ccX8JW4rZZTVqfziEHelOtkS3B9K/pW1Ba61wF+quhzv5ynC10j2UNS9a0hv89lNEy9
mah/CeZa2X0QogyJAIfI0qN3XuPXIepJBezISnwJm3p2BkBRIkrwlHPmvJpWxM7ecXAoJwH+xd4I
SwredqcdB9GzWpLSqvdYv7xRlMAsMKDFNO2LQLvv+JCBE5fvzFOEa3rU2ScTvLyof/GCVlJ9MI4Y
XZ8++UVxoEBEgNhL4djV8tRRfwhOACI8DpBZENHr8BORdMe3dnRMwmlb1ANzpWBUTAU0YGN5oGkI
CxQ7dkFBZp6xIl/3ca8Wj40yKMjUyMi21k9p3AjFInkg9lfp9XIpqpdUmrMdSJ68rt7trIuBAlEr
u/3/Oqay/o4hCd1qRJ6dPd67rvq7e3dBQcKum8aiY6Gmk0QYc30x153gSfpEyezjxWqBMBw7yvXh
QI9VfyDekK/LCyvH8IfCCtwQ2aUaiGXnh2RwRg2sirUVNrduSJQsPw2OkGeY9Tq1IWY4ZelCxEgN
THcB4Q3VQL031XCjkdzAaGSxO7+Xf/ZMiydAiapz2ekA/3DgNyjLTgwTdWWyTh48zZ4x0Oa/yWCz
ysjKALqPY5oFmReVU7Zy/rh9fmoKw+IjPRQnRqbpVgFONlhwsYeHUbdpiunOnP5c3tHhIQnMqwR8
lRH8BmQhZYzfVyjotpGUUPbJYGswIV533bBIQXXFczQ0PYRKedpfu3+glgS6MziJQXOiCcLJoHOL
N2kykvdG2TsCEoHSKo9qQhxhz5ayTvsLIhHCq29u5c2FGIgTLWcLOYloQrNeBX99i9UmWcUZpTIS
hoLB60ySMxMIUsfxZmZRBpfVOQ9AKUMS0/Nn4ww9qhtVoCxpIX8TKOjkqA3JNw23J3ZkxUabc4Qi
9aPXl2X1VNXB7Wh94Y3rO0I/FThw2Ut3wikNoTxw3UtiUMnKpq8QqloIsdUJ0MDjp9SZLVW9qsdK
+TPw4IDdYazvpG+oyKiFfMlP8bvOHnyEeux6LiacFx7TlzojDqgCNusvmkfboW81kARKTMX/7BMe
snNjlQ54iSBpVOXf7RHcbQ06LqXOE3ulBB+llbwLA7DEnlFMO08Z0WIdzgIAxYuFzWOovsf9kZMr
AIAptIMM8o//qW+F7OkVAe6BXJElr7pgy8hVw0GSbuR/dn9TGo2CxahNIfiuDY5xNFmrPD5VFX5O
PuIB+3UdbdJ4ld95+7QGbu4DPLt9z5XE+JRG0kdGojDD366rLQTPXYEfPr72X4PU/fIVtnLZnGEH
Mhn3My9TY2GNt+NZV49q+xVwgP6jQxk+nMcQEpGy2N7P8G36XYoobzqox6MVbP+CvLbKcKAdouJz
09bQcjbpKVWvfpIFCebhzGXBZdKKjNddrHxlR4asBPlv1k+PLnbKW5HHtYRigNNlNr+9SsBtu++c
92b5x/sFn1LHZuwW2LgIo5gTs3RF/A7SJNTqUSG/me6ynsv7QSp0bUq1/rK7p1Ctw5dXOeKnsLN8
jaULJciAE0FcXMOXRbR1vUEoJxloUCvsuRYWK7riEUmD1NpkBd6yxEblpWZZ6uODS90ilOd9jbSc
cwYHC/PaxT/pfm8UlY+HSZIk0sk52IPMzsU19aXaDkQi20If991nEWxJTRrUdcY0zjJRF7OppVF8
eKtz0sYx/EP/RoaEOCxJMwKjL9X1rBXhBSM/+Z97BFIUn9lgl3+pwF1ci9YEPb1EWtx+MH0yurcr
l6hty0r4mZtkqnsIZ0oCHZ4yJsivDQUoyQdZ75asILEING4PjnEG/vykhpw2KjDv3qccC7UKkuQ7
LSMVxDNmEZzLm5+OZY0cge94ohOyO7fE93eO9QbRpP5qc0Mu8sruTU/YxYx95RwMRChNeKQLulbC
dHuP2BZSuuCSQZpxI/2hNtPNiRBM1apbIiLwpQXhlHZWca4IV0sYJEa0o8e4EMOjLCclzCePNa6E
DP3t+vf8bzcmJ0MrIQw6H5N2q9m9xJ0IDFUueoTENRdDQK5Adb3MprTqgj2dtWOdDiALDI4zPq4k
nJdBDMA5Kqt0CE4re500CMfi4HjHMf6HNGj4H9Yt7UchXQJnqqQNeo0oUheP4VIBImGDjy5AwiQv
6yTVDNjslz+cAVMZ7La5sPf7HfmH+I20eat987oaiOyK8Y+yMM/dpa2jEL4Y7pc4uUeE0N43+UxB
46mrogBT3RfOfyeFwoljMG+P3ysNQhtMDI9UpAy2VSf/CNDc6RO23yd2Q7K9p543+mkb8Fs9E8Ov
o9wARfdHd9a/b5H3vS39lC0v2SGnXT6sWlb2UQ2NyHYJVqD75ba57VBKZSUMqy8Bz/Vu32cDRoKg
oOnNImYMDDHYJkjxfp10WLEjQ0x3m+l2jb2I+GdZ5mJgurfqU2Er2XJfsTF1VBjfayWQ4jTz4FHf
3+UXKQSRPY54zwf78JjGjCPgkFUmKESzVrmjMKXTWyV/AmfurNvHMuVrsdgusv5S3nSJ+1aIJwYO
fmlKnROndobc88LKe9fdGLuzovE0zdzqqJJRqFDOXP8It00klW4KJy5cGiOjLjycDef59MXVtSTo
fNI520krih4zlPFZHNnx6ZC+XWPLHLY++H+dk9Z+ZWz4QtI8oQCYysa80EIm89uczyr39JEeCG8F
PFuVGbMDX3WciSRLi0O9P+GWOfPz+m7o1qEkrwvLiGvbbRxp79Vinx7ebcild5dcJ5IRMaoi4vDg
hO7ovTYjIrJVpDkL5HH7EZm9TSj3LfiW/eGhieLsVChYx2y44+NyIZzEXvjUVuig4nA2I9gCx/QA
Kz4MGSwf8IIPDJJchKz9rHDfBFSZxclu2/QJRUeP8QyCIHAMsbf0ja1lXmu3WbgQKF1ie5Jztt9I
UgdedzfnBkv6ndiHlM6Q24a0/U5fBcXegfIRmLlmvO2U4cIMPNxP1xbs+LTCRkH/GDo5TK3UNsUL
fqgG38nQYJB/XHfqGheYj2WWO4QEmTH+ezbWuoWOF/DG8q+2EJFG+tzAXzY1ANWfyaZ/6xXWSpXa
fhphOX2gpygmGxsY/YapwtnekvDuVzJA69+Ty2B0oFUelGpmnSXh4blMBZTKK56nh2XoqNOhnIy3
AulMnGf0pSYIyFAaeEfICoDpD9/wmpEPzhTXi9hhJZHPsrzt9FLG8XTAY8XXHetDIsoT5yrVjrmd
l59jZfuw2JlHKEnH/Uk9kzIMz/hc2NDudnH9Q5t19Dy0V9cPkfBaoXtvK+MprBZCGkTVcRWioFKz
i6ALRzMkDbOb+pHXgcpKN9JTi3k/NAnVuy4k6IAN5cQpze9Nl1UvzJgccKH2BkzVtwaFHWspDWSP
S17cc+BO/DoWOU7Xbn7fnvFbIUAx2tLBPdDn6cxVctWcZOqv1/boi/e0VaNADdjKnIKIwpq70vhC
cHIjetwZfji0QyiYcRVuTPiSC0/v6uVGxt8TkU6ucsKkPLrrrhMTYTnkID6df8CrciOI1kkzLq0j
cWlKYEt+BnTIxAVM86N5NZFEdDTiY40xsF0Caqshc2qjlz9bc90xi9DqIRmfaJzBI3ZbD5UWBKPV
yBChRNYNpMPeiV12XErcpZ+BGAA3mm6UI7KgYtijSiMN9XR9abLdU1OG0qBPB8IVRXxLtDDtIL8/
qJmUS5kh69lzRYMY6DfNVDbzZtS1I/EKniAKO1HinvR68dNcEsZBnxN5J28etuqmzFoFXz/u3s9+
JDWfUDaUeEqRTdXniXrETU+4tGSiW2tnUKNKHbemp0sSmhcYZWveG0LXUPE51fFsnurX0oNjWR27
FvqdSVFIz9jDMEmNzMx6u7oHFYv8dBsmULTmRTT6kBwQVytwHOkCmQLjWn07A87pOFCSefKNGiXl
K9EigFHkdzibTUQOogn8vz5PH+jNDo/H8VIv1alXeIz3FtMhgiPlPwc14w3DRxwW6TDc7D+KfsK2
tjPJrh1qEsJn8I66pnzOo0rfS7xYFgc2NrJzQYwHvWYlFS0DrQ2W5CcMJ0WkH8uxLCbCjW9PZf0R
7qKBWZ78F9bppMonUb7mYwi5+hcrNxIeuu59m6kmmr7lXMsKSX73tdqeVb1ysV3eIKh7ZMLzOGwj
d0walXOOzU3/0DjceN3N8LIWhvMyvjsxIVs1SMThuGpBlUqrVS+B6pFrdqqFC9DRU4YbLltbqy7C
atQ7jBoylDVRruHUGPI97VO9WtgAI28jdhjpiR4N8nHQsSgdbW0NEzVVwk1TaBv38T7mUX23eOjU
g6iFVkXhqf4sCDzVHSs2eY9EFmWEjXGyNdUNyvFgdu3NKWrVRUpYqEHoIGXgzVo4f8pm1BpxpW1g
1DDn0gyDtbvKACm717z4QdvjjcxGMDJitDn4iJOaXc5isNOsvPTGahuzIDporgSXjtmk84nV0Qa8
gKPSp3XeupgyCMG7QfJ6bOskWhJ9HRf14nJ6xfhEp3U5F/x6OpZGtJb00RDLK5HQ9Jl0k48IjBgY
5ElhhT0RlugnnLbdZlzdJife+2rM+U1kG/YnZOrU0IcehViByp8oZRF4mBRuqKo6oQmstl5ZSP/a
KgSWpmRfQVrCVJ1+4Hu/cZhsgD910W3zIoXDcNQfhh75TyMkr2bcRIwQCDPP6KzvOqoRDoP+Rbnv
WAN0wbgttId7B7f6i0UM8hafvXmura+t5X1mak5wF+lG5kYeBKP6p/p9OvGteQkAq/UfwFI61s47
dKNXqJf2x+LtlUzKV4AijUSQPqyPRz8RZ5QxsI4EcJX41jUwumFnxsGTJSr+XX71qgvq/8+sc1Wn
DTbU/tma1K5RcxKa9OnBcT3KLb6TxFzoNg12AwY/0kh5/McZVL0VJLMlt4FOqZSV2JGVXWDUVVDr
vl/os+Un0wE8LTE7EVd6HlVYxwk0LMon1OhtnKkRg0lpjTRErmbXc6MOOCLqROchuafvEwPuVDL6
3Jc0Y++yAPzpomcjNvfz9rRZVlmaH+ufvkjOga9R1Dwfh6CNLOqhMfPRmuKur7r/CPBERGyPTNv5
kAfzG+Ks43+faqd5J10qCuzwRCjn2Sx8s6PQmde/byfS6IS1MTHq9zEpp8lJRs+ktXWko5sb9j/h
w/PkU6AbVIRf9UIRM91cWh7rNxysPzeAH7ynAD0Zb/FjcmImbwUR1PTgtQIppPs9c5JzHTJkB9Ro
GR9+IwiqOJfiGtTCakj0M8uSoG9s1voG1p0pYlDS4+PseX94vtOvl0glbuHAdRePJmjG9iwTx5ah
8P0/IFADkL9LcEKAuJ92wn4287QMi+ZkRVeqypTcCg6smCgr4XtCV9TJn8K+KcsRW6F+YZh/UXXn
Q+m5vGAeaNI4R0jSMwT4f054smlF/ZPBcBh6DbCDLTgPYQpkKxXGqYRNq8ZmNx9f9LyytnkhKo4w
RBQH+oyaWRX2ixVbtSHSuyN3b1FaO1c7ornXS1pppuGvuXInLtUTKw5DQs+r4x0116w+JxzRfG5+
tsdaTaJIpMTMyvkbYrMZhQ9K2ZfSkzWKuiqWkCPFPkA/0os/zVGZwBbXuYVRHgtG9+zgVSc3mvn1
J2bQ/tm8Bx1qn7jIvB3ajHjMlJSp+H8k5EvB/Hws66kAhXdIcV+8W1cewaspqZP8i+y2+9tSxoIu
bITRa2zAVsy96UHpJjjGH/r2dAS4XjpQm42+njwBYKruQRpGLnCspudgBXIRISxZ1kaOSkfm9/+Y
wAMnxzYaigs5d6dn7E63Uz2XFGx+RaUT7KwdmaPaq3opijQKJXKsFDQCdx53l/jiJmgeoepE1uuI
ptH+HoEnluMj72RUSlfJGRpZdbkcsO5gYhJM2blLt+NgnQ/Sb53dIH70zmIOThlYEPVMAdy80ypl
7vNz6lPyg+HCsSbN97zSWSWMBZrbnBDIbAW/wfuWCC5n+hyOZ+xrwoGMIT3ODtB/7KgPjguHw/Pk
wgau1/v17NpzrtmIcacz4srlLh0Jhoxyd9gvH6M+Ay5PUMBSJg1Aj9AKjGMTcQrP3jU873q2gP3S
9iaOu5/Im0C7uTrk0mNxyI7XDpZM0dFwbcbhHdeZgVH1xmbUlsZ1UuR8XsrW/oPpfJHTaDj/E7Od
sBsYJYTNZFTmZ3w+EZ9i1kRox6NEJnTDEdKb8g/mlBTpRDD5sYQZVoqaLI6KNQczDlp34uwlnElt
Joh8wmrlbG5wD8a8Jpd3mPTOdM03KFzv6l2OSZs1L3CxGZnSxqPmpXFmRv+5w8wD4XnXYCwQR6pa
Q6Pa/OjIPTMfixXvSBiexHTv5AFU7ClmrqWi4L63UYgxdSR3YSYWV2u7M+hLktpkTOAO9edKTuei
eRyOcjvUmjlFhYSnj+7ewFdHm5spgNAol5r2H58tkX7OLMzw03AQwfxudO2goJlc9+LAsp8UTdKs
+7yEZKXlhlyWj4Tv/7DYwjfJn332JSGXVdiMfaRP1pGb7tn0qcwA7sbam+JiPzoBoNgMdB68L0/R
JJ3uM9t0yXAnCrpbGr800lpeYb2Ri84z9X0zT3rEppD9A6PWoH2tTzfFUj2Y4MhcPmom4FzJ038v
yE4C+Ysr7gzc3Vi71H5Fb23we6F8eXY5y1AOD9fiXzWBaLIbCVdH6/TlPv37oPMAU8+IponLXttd
FbasMCHA4U/z2kwiH8jr9wOmIb0D5E+ZTx33x8+eTS04XdV5buxAy2Td7q3LVzmya8oAdF+kjDkp
L6GgDib81msfLEuaENMmOMRAASV5MkDIScWwAUdELz23yJcuWKIhw0vvWk44SbFi3F4uFGdqeTXF
iI/LZVeHMTsjNe6EbXED6IbuEhn1l1o6pUBQZHfbEZsE0BkKN1n/WkvRY/EvXvkGFmoBWN1573HB
2SLSFBHusJmII01LpSIQAgkFUUzVUTH8CqYDpNBaN3Mi0XErnS+7COW9IC3aSb89htjCqFEc1JXE
A90P880j3Metwm7Ps61dcjWgAfQk8EWmxuUucQcSXN9sN9IR3ycCLPlbOF1FICOgZTWReS7e+tJo
7xERjMA8P3Vu8DyNRSxr9pYX+Q1IH/RkCQz+Rpv5lzq59q+e5fofrgxvzoBAPRygM/hyI7pgfISx
bN51h6w8V1OupqXkPpVptEfwY9kDSi+8lkd3CaLHC69m45aD1OnAXdetIlUzd1nRAeRyQSmCBgEY
1tCqXLhFmvWS2MKSffnswaByrg8Ne7YhZBuMW+N0S++8JFsc5HJAJScO0y45OBU2ycKJiijcwSF1
5+XN6wHz6sqMW67vRZ83bbcz2VkJBO2JpzjYNbppf96AiTM5r1LjSMER65lofJbNt1QeLrb8EInP
LZnpkWiPNEX0b4zRbJSG/27zA7qW28m5dDggZa05PVxNMy2QWxJGqU+MRDfQbnLmcRt8lswy3fS5
3A/0tBA6rSJmGbGYxSAOmHXykZMYRjDfWIwzGlQmytwaE1F2LQ0SNMOEsX/RVjB0x2g/sF/wpYb4
HsXLE5grIvq5/3YatdcHeWPBaoMkvXUX6rYhMUKL5p1raI8Xx6Q0XyhwmBUCZo48G0tq6tGDCgPT
yJwFgAOsoTO2JcP/bNF8VavOGfhJo3kBmvbnvmwtkBXnYZFWymVcFWX0/aPXPXDSWyBRnlsrH1kf
bcvIfOV/RWUtDRVz+ch9dZPv7l4exqDH+DIdIjOJ1oGxekFRUdoNl/hez9Ht93iIli2F6lCTqe24
5QLfJHNMd1lUNqxgWT6J4BZEVBFi33dCE5m3DPvb5viRgdwwSNTeaUw290oeXnuIdJFJjtlmbIqD
LFPgdOfJbecidAXvwwT4kjg12YlrT5wmsWqE9NXqRBSGSV7KBzp/sCUCvsMbmr9gS2aI0JK8D+jA
1L6A1Zds+k4f3pmkMJtObEZO7LERMo+W15j21ujSmUP214GxGiRY0IMJLhaX92RhNrduVGC4X4uo
XIXSdxpmtDUYA/9hscCplPFxpdy9/ocyAGn9sMDwajdR95pFPFGqM7rHw5UUopAsdu+nPGeetCj2
33DVvgBhukmvdE9aULJP8rwC4WDgOGTu4TCeRoJVFJc+K7DArn4owaq6S0J+Afi7War77Zw9zfoy
GlFiCdNG96yh5iATAWcxHZxwq/4nAInx7HfcW1+vKxv554iB/88g+aJsxG7mqrPpMHH/wN/X1AAV
ax6nTsiPljwUnuO1gG9eEo1EzB+wcaZr+aaMnTRN7xdSsm3vM3lKxGcclic47L3jfJoYsuL/yRgT
Jyt/ilepfvLYnmrZyXY3rBzWzkL8yw8calClvhHNi5+/6AVtg+Ek7Hw28Z1cAwW64lCBOI5RfU7+
VglxeeuhLOhbQnS433LpRvqV8+7Y09sHA5MbUH9ovYlmJWIRjLWokOEKAjZ0gBt3WuRa6xatdbm5
WXjX5h41X6k0ziCW587LmDyPeAMxgtXbJzphqoB9+dP+dE9CQtbh98Q2rxJ6ESifJ8d5FjRY1qTq
vVQpXID9mgfrxVBPkeoHyS5+/utkphnLCP8LS3Q4jWObXezblZNYbzuENKCTJUe2QudwGPw5LcIj
v/n5Iv5pxK61dRJUOtJKRDE2X24IxaUhImN6B2xv0eY3+Ja3l1K9Niklfmg7YhhBz+NfQislA7be
PGhpkkhcPqUpxjRf4DDa3FWuP09Zf88xINovAEHuZe4EfOJUP3Mt27Qh4wyPH7p3ZA29PJmz0mub
NTY8I37MKRQgoeqvH6+OXr46Jqnq312QIevcM1buLHiIFfQSWTMMf5dMBhpr6G0fk32b0Xnq9/Hh
HZHSdhSFleZA3jjYoRrR0DSIf0P6341q1v+2Qf+pISGcyttAOGRPYtaZiX50Up/GClWfGKXYtMLo
ev/cL8BdpQv+P2hQc39X0sIlhJ1NCTgr+8Ha6sKO37JSDBz9vEQUFBIdbfcxeQ6yD+yz+YTD7Jvx
BCEBzyKbWcLUOiO/x/e7C/xVjOwhrZLUZh5WcF2PdN1pBoPf6v8dfiYCBDuvJZDjynBfOHHCezec
T1ww7GQLqaajRM4nSpav8Y/Q2JT44mmHSOnb5ogcRTyS6mFqe9cUupJeHIzMjKtrqJh2pL6KGA5E
lXsjSfI6jnh08YCBf8uhmGr2hx9RxhDPCZ1B/giG5YsB+tHXIhE8lqRoiqxiK24ivH90ECfGVWM9
TfMzVfir/fZk8cm4rNDSxO4Ezc/eVP68s1f4rYPyOrPRagK4WeP54XehNGPTbAyPPhDLHBmeUAcW
h3H8Ynh/OItdi7nRYlxH/BOMoJ0u6uDW2kyz3SZMru5aFNR8Ru6MKME1LnbpsE6lYZwGr7L++MLT
NrAyVPhxPt10C9IeImNC7OiGSToqiFYHxRFz8rDGWP/PPc+4Lpl+jQhYcGVOpw5wtv5Q48q7ljEW
peVzqRrNTf93/nHnJ1jM/OF2aXDNZVEX+uZwJWc6VPzyKI/mchrN8igIqYMTGZyzf1m3N3A1a54H
oPwDX90pswIEDry4+GPvsa/0I2FLBcdFsofeIY+Jz7O620b+M9zJC9xacJvpGidAaWnM7kszcrWB
XKff9IBA69TWmpFA9PNfshv8A59tEyC+vVN044YO6csJSRSGkgDVrOWbNtws0nTAy+YaoexcSyfq
zB78L1LW4qePu6np5ciue2fXqV75TjR3nPDJwz0xAwt7uZCmjXKe5T6Iug0PP0yA1r88+k5jB/vQ
VmsNdELuvzt5/jl3MWVDhYQrElGHvtreD5enLM0mAP/j7T3kr9nvuzdUm4Ke8VniVLxprzy0ghqP
QHWfeGmluJLT5SjRdIRswGFie4hWOiLazDACSu76LY+U8S3ChskBZIwGsIZSOdrwnE0nVtPdYWMu
aHjgF1XYD3DZ3XPfz3ZUI9qJFOkn+tU7bW1Hitb3jQAEQG4vCWghviTHFH/381dNTzGVcFGV4trL
QqJyQVHKzq03nchwsNgxVq1bf3ISaZHgJl1k4Hszhs7HRKbbzW37ZGZ7CIhixuMxT2VST+yrv2zq
68fS108bjIbhA6BLbKYOCX0V9tYzs7o7KruTYugFHQDiYU6EFs0bv12B85o0Kxq/RGuujAsnm/xh
tGne5PvVYfGMYl4k/GxvSnxLPo/J9NJdQ8iwFd6jHycEbgaCIrkLs+5zPzWW0yfFcCS4Jw9PleGp
fQYhPaHB+3MgG4H6Y7UVzoFmAvUNpxA6PY+XXehvRscnKXt+VA6HfWTO1vE09RRCnztOziejDs3j
OLSrMC/cR2uscWoS3Cn+OZcfmlWWTK0cxxQGa3IjyN1Jry9UAPXJRjaxFnn7KcZh+SCRpBLT4FpV
YJYaApdVd8oU3F46BHufNXPWhyDcwYbxKdiuTk6jEynBbqRE3ILDAzHhsRIF+mkrY+i9BlBMkVHK
FZHvJL0k/JyK0EnYiCBOL6UC77PsyJCnj9eaF2qpG8fqPmmyGLHPLDjoi6KHK/68RpvPwIeiBcq5
iAozwT3nHp7BoaMoHLwtRUa5tHbrwQ5nVIIMqhwp25c1FxuIEZKZ+qjBVlpTuBYPN4nf8duS1o03
3Nzv1SIUQl0xuldjgBxzkQa3AMturET1+3ibxWUZ7GZGB0Kxv4JAtFWiUWyBRPuwSggTBRXJyf78
3Gd/YDuNG6xqo05uHDMvEYqE1FS4MQqKVpSw+nLaNzyh/c8owJfYYFagrjRmeFy+S4YAMGYG9JfB
IPcc7oWoBivFDsllNr1MMEnwe/qwMAq8VKh9V2qRPkAsw0keUABinAD0gSEbfbUxZ4RMd8keB2ym
ImiNrPngJgXU7ubywBB5R2RCZGVuzkPXlkpKXqr86H9HZbBCL53Y4hu4HwVnpgT9suYk4Zk+9Hwi
T0iHViu+Wpdi/lPL1jqWRJTaz7bsoINudA6geEksu4OjVVhHGSmKbOIACf9B9G043WVEt6MYxIi9
UwWgR0zBg2ywoxbhzZgBf+E5DBV3rv7KK5YmkNd6B9EbPUeqjpWFzIi2s1rZ9/36fFICW1vlLNbu
rD4JrayGm3kFJG/MhlLtX71lKc879eCiWDfBd3GtGGNHWQn44PAKuPiYvwFize/lUrk2XxDrrOjG
kSEBew7wAF/Z4XDwvCjj1rdkQcO+9rRvusOSbK3CIMUXlLY5cm+3K2TGb8ezF5OBEACPyw1R2RM/
FqjPilfwXi32HLYZUSkgfnz52TZCZTtRGIkf3/M44Taed60QsGe4aX6WEpLPfiAhUxdOClJXiAMp
tlluPgTVkh7Eos39uVGK+8aHKu4+UB4YRoLTmjncub7DgiKOwcI/nwPEdCiHo06cNVUDDW3OSJYA
oStAai8b68fw1SudyKEoFeH2Mu+wFqOmFtPpkSCian8eehTkwHWfyhs3xh0800/vDppl7DazhZd8
okRHHzQ/2QJgQjieuGS6zQK4WQYWKRJPIWyHpr3Q2vsyrPmvshqx6m6092lvODvtU20ACj+5stBD
hBN+P6hyo8nT3mq7JGBQ3zTVf89LZv7z6/EH3LI1f6sCroL+BmY5oOeeeFlElvQWQurg6Coju8eO
tw/DpEcj6Th9QxN7hE1JLZwQjDGi6PT4S2EYvw2tFwEKF1peBc1KpPNZyPBz6Jg0pAz8wVi1CsBG
9KaoylIJtFMLQwzreHkC2YTnhoy91liCWs/BzvWKXtHJO3SxPzICfUFhpXmE3xwS0aFpqlz6qpBq
mV86bDltkJb3eJkJMQ6TFxbBKVqv7djiJgUd1Q4IGOkdXZ09o1pg2p2hh72PzXbAmKLq2N5jANwE
L1l3Cz2b4lpXLHB0aetUEBpivYNjmawHLA65JwGaICNmYthA1iPhmVY7WEgzRmEU+r7s/E26re8g
RsF/whgkO5qt3XlEPi0F+bWjF1G51fDgi/sXW2AcSvni2ANAmY7xlTMHWBuxPjCiJR7qh/7Qo35B
ikUSEM15af8RYUHsozxkW7gEoMLzqHUWgmYjPhnMg1IBERC2xQ8ntptvULKidt+qsYIlvU5RQGuC
ZgOkRRXHXagdenGPH7yDkSvRTzPZgvFhGAAH2VXIaerE11TB7BUIoz7E7xA08F2YM5cpb1Eq0wf0
5jzeJul051nFMAjYRZOslTK/5O0OdkMxnEVueaZX+rnMaBsZyiSQlEWjiMa5G8jaAK/GmYz4qMvi
8c6abIG1Kq9G8DaA1vdg8C1INNvBnA7mIQs/rVC6twNOmuPxN2xM95h5jqGnui7w1ERVQdMpeF9A
QNLyOjqj2nSlP0qBXmTz7H2a95t8G+xxBj/Z3RbZHXcQyycPb09E+ujYVJuMNA0V/g1PRbdegp3E
yIKCMojesjBbbc5NWpM453bvSkphFoHCRhqyVbzMQNeuNKOg9ycA2Wp0c23OlkwyrKPFZkw6Cvu4
0ouJSvgeNfW0xaobadr3iQH9t4wts/dlmo6qSPQbfk1TFg141/wZVrhnwNah8s+73U/oYfqenvZR
8WXfMmzCo4VGhpxaPr/PdPO6e8QFUCl82VjLZjzwP0rMspj4ZBkXBEO4fmDpaA7c4hXj/aPueefL
yQF6HP1TKs3faAcuaXkmvnHJAKhvdjqxzDQ8Zq/58X6Lfc04hp8GwRBWCd4z/KDkQ+bowWrO5y2T
S35aPfroDCrcg9lgYa/4IIELzNTdfzAXvAuRSsy2AujnaiPmpWeF7PQpJq6ar336O0kFJAL4WQ7L
WTVQ7Oaspl8dbVgntAkjynkOG61bDqXBpQQrvG/Qa2RfCexO6savk/aeZeFpMe7GLnY3G7ebOQhu
+872XNdN5YXi9OMgzeDscsXm2ixS8fVrg6mfp73c/LT3pEM+kFgp/aGiXdiFJ2AJ9zD1fn1k/3Go
bRBUN1AzK5nNnWjCMi/5JwP2/a8ERuM3gEV2+FcVx5Jh8GDvu3mKicZVeunWj/rEc5gdhnmLyOkN
QQ8SzIrSFZqwSa+ZmTSIgXbPYiQskUOxCRZWp4JeQ/zI7tbXqfRrJ4vevr6Jv5Og9wEjYSyOMhJv
5uwWhm8MegStYlt2Ki06H3fydfcFcHGSKvlxc+0iBM7lxf26vMeGOiOu3r8Wvmp/RYw4p7+iRG3d
7e1JJm/MLTjZlyEDNK1FKL6TqaA6jY07UOfb1jCANu5UjSyZsrRQXWZKnceqLo4aeHRELGOS4/Q9
V2jM0TiuPHZbsrCWByhuSDUHeZykI/nLBDslvJb6NSxlx6V4cIi0guEvJG6Ibp+ouWmt+0Tbiz9R
YyL6RdwWMnRaPGP45MqniCbYjKb3N3gBJuOBac+ywiXlGhNNxLLoqmczhQVT0mCzuFSYehHQIcvW
pSTppzkbkaaGjS1iDbCOZILTR4UKeB5KE7ZE5nzv6EkiREJuD581p+j92GBdBsr1MV7rqscAZK/E
aph3dg2KE48kQYJsROvs9v7tSJTjdHGBSvqU2CU7iov/OPnT2XVzllUsyBnxc0kYluqHnHBFRLRO
5rRdaRC9ezn+vnL1vtROgs6ua6B004dkfXSkrLOiiyiQB17oTofZ5KIXJNgjw7/wjXN/m0Y/z2K9
Cp6gqetiUwZolmSk8CteMLv7B4cb7VtPBPZTqWAr+sgZ4ESRGObXICvImlXX5PI1CEL163SsEX1R
dQtjcVrhN7+V3BwAelFL76bodK4qWEG96tyuJTPq5mOsCO/Y4MRijrr98CH2jqD/f0pfMjI1iV8z
DkDLu0DdDLiYy145b79MRdjFFRSdrQ1ti2WKb5K78sZG6YTAaqTMgMbzn3t1rU/a3aSWUiZssZ2B
iAgzOKVekoPBVclTsAd22Izoa6j1eUPIEK71zURXzHHEYSC2ovYyJ9cJHAwDxQAyDHJmlyQc3H+8
sE6riuVRyvHtvRmUqJVXH9oBtB6oq/P5pVIJtrUTd3ndF4MiWz6rD5CIq4XTzFkaBBBSzSZELULO
z1lIQ+TEHF7OM4a70ceAt+ipFqYahKqfj6eqigBqLwRsLWw1K089S3m+6qbM3/XyVfowcU5GzX/c
Xe1i/W9rr8SlJTPdFrs25fM+oVZ8J/LZ+hwj9ygOyrBMxqEkoIpUOLuxs7kvwy1Lne2moae3fk1t
gWOzCiIoKRhJKYx1emXN6PyTiVt17Ce+G8+FMxBGOJsPkS1brzTpE8Vbu7bjmnE4TOHgavSISDri
XLzxx3fpb3+9FYZX46FiGTS/Ka1RkU85Y2wKvcgh8Y6QJ0+hI0aLdnFOkQEGd9FwQxA6LgNndufv
dxF5BPo7p06lHgjZr5I6Ah/g5Ky6dT+/lgAr8oP0DhUkMxsqcr3WuvQJVQN7Ltb9IRw91sAkstgI
CF8R1GHE9bzJvljLZA35s3+UnsVIj2sWhZyYpJWwK8UGQCkMpkXJMJBsJVlAiBBY3/oARgcg7Y/r
D6ErB6Bz1wEG5sUfHuSvRfCMuCaCaf5vNZh4XLhYSwfJLbaGldX448KniE0EVqN02NdWU7eNj+iZ
DBhUjuravopyYXU9MgJeRp8tVzi6AGtdzN2MrQV4/4qDg/f8+IRb89zW3cs8TVyFGe/kW29gto8v
Bnqid1X37vL9bSA3oxd8OF+30gBy8qrxd3i2iTLkUjz8UqKgK3AqlFukrdLs+Ue5YvSfsccmRfpT
dth7oOnvEc4CjNOXJslStD3VXAPxVQFdodf2TfS5i2vcefwQg/EwSbzPXELXHNpjYtWla5ApvHb0
ikJonKExqAS/A2EbuyW3pHjEuthFM1Uo7vnBeUItyOlcFhEMV8sOTom7dKr6ZGXgsKIfSDH25woZ
1Kytnmk4oSapSwoBAAHwINhtdpUF3QQ7NxBFe0+Nak2vXhhXceOyxDfsY2ncJfoLf+S5eMenHZLj
e9+qkCmfwuUB4ZKoecRryEtHI3GWUexpYKadiTCPh8WvgE0Dg6XroyO50msOtNsAQvBvFHgpD+HR
OixODohHfrDs2IsRSuNFptrw+KT2d/WBJQOU9hbDjEjYAjoldy7cYxqzR/TQDsQlBPT7stBT67fU
oOha3S2e1hiesivHgFtYj8AFPkdPaAJ248/Za2las05xzgFKflA+k0R+pOK0XE0Lom0O9dufYdC6
R3jk2znjfb54sAv05LT59+CpNj6YEZvqtFzze/x6/qEe7v/O7AYQN4e9hXscp4sPT/F1zIqgBEPE
0YxSgHEOTLqm9YjZU6W+lY697Oykn85g0uIvvZUW+EumHsVE5HOvwSRnEtwT7nkzhLVqa6QQTBwH
it5W/SJWJVv/7Oz8lHEx/G+ZSsoQdE+NNskuwyEy1uA1aoTmaxqaDVZ8rHSbUDaOPk8vNn+iMaCc
oR4glIul8+KWzsxm7XdjxD/tFYVqPvbQuZCAdpmrRGlJP1AraIe23CJkN/FVkifLRD9cWTPK0+H9
uTwfQyl8WL6KQv6kAFi0wOb6ewx6AvmdTPJ/m+ayotf3oK8RxjqqMZ5LPR7o28AH6D6P9X4pnzy6
PeARx8IjWmBD9n1kfkdfXATyjHsz3vuHftiI56r6jczIr/qXywj2jfDgl65jaUwB556uf1jRAfEm
d+sJ/2vM40WMSqWEv2iMLq/VfFy9tbQfprCGm9jBg+lXwAoNi169XZSk9SC6M1KcutoB64TWVn/y
hMFdwxWfGGQinCSZ75RLe+/GVoNc6nlC4UC6b2rhLm31iUEqaWz3EnF90vV0rI2Q2rJQHH3pIh3T
39SAWDk/ndvrhV4IFS4A3/ohNZNkeJGYsQ/B9yRdsJNFH003tjUbLZoqTR0hKR1NSiejnTvlKy65
Tux+c5ulCPIni7mueY8xpNfg3LfleB7fJsoisCkod14/GoVjkzdTp/RMxQPzfFkyf2uyKFEyEYic
BMfmk51X/xh9nWYZYaTaHBEJjJ96+HZJmg9RPP4QfKunI5btbjMPW6X2mms/1549lF+uWIJSfO9W
7K1M5PoDXBPQL9OfH+OZp6IlWez9JrWm9IkxhWr/2hVkZk4CelawhOoYNCNkFMCWCURw4Vt3qSwT
/x+HXZ80EHjJsi+mIze3RX/ffwOeFioxNyFp/OsddB6MRtCzG/pwYtw9YtVQ43nGNwx/osmX41Wq
gj3VqatOetJZ2Uo3y7HusgiZug3/CxXP1nur0MFndMkwLIJyPWtaVrSw0AwGQVHf4hthnGY3rT1U
5xBe02eNrCNlbszpvbCjMs60RO8Hf1e+HbkUN57n2j0eEFORJJUG6XHWLVwIpG+C0fPMLh1fxoiZ
PmUn6mMOSzcqmf7eugExszKGt0xca68vIO+/R1LFnWL5UgJMa3P5nGmBn22uL1ReuBzn1UAoep4R
B5doYIxHrt4nTB7e+bVREoZtvL7NR+EZIZzw0nj9OYP4JJhk0c2v89utyUfvCydu5TU9qSyTaJEL
qHGq4hZ5dYO9cwMjiS4Pg7Fs6SSIXXgeLHzbriDMXFb3UfHCLoUZgp/wd9wk/Rkdp8uXTHzEFUMT
bGqKQUnmyDlbvtwKs68v63ClNlmTHXQppTu2TN1t9RpNQeGg7vgAUus4jKPZBiVND1TTYaOIEgOI
fHBTT1br/HZGyi2qFv+dNU/aYrZ6hH9m97rLBC55QakFcNcUyBQzR+4+8f35GYvCoRUiIah//NYH
9Pt8d9gzia2ierroxus76gOCLWW45zWyWMHWi4teqYVlAPIqojTcoGihUuLYqYATOe0AWQcofAo4
iTtaGCM8bLW6Md2nZoVlCNLdPp56HbFiImlzG51Xjc7yy2YjAU78URaCIt4pJPyViTGYsHF49j8r
1Uiz3QuDDa7BY7mE0ez+bTRIunexOOX5nPzbyQ8Dq222i/QAFL1RyqRtRHsyg+kCsM2IYQN19VLG
R4tAW0BeTIco3SjQRNtn6C2PGks7MZBkdjRQZqe6n0i44C2AsewRQspQ8kwYS0H71/SuwBY+81vV
KY9nGaWykDwc94/RYK0N7Tqr53Kk2ZCuAseNDXcVfn4TIjU7wLzrId+E2XvhjtJabZzqc4RLxYxg
fzJ4HT1JT20o0CWdmAnODMx18DF0yq4FF6Xieri1FNix3BdRTJ1tnjmPAFzcCAghPlpF/5rERT6h
9ji8iXS8IKhquebto/LUvPSGhGNVN+wxL04Vu4TRkGI4gwc/DJgZIUtuY5OvyKQziD4uR+651IaM
ziMBIxiDrbuObdKyMPBh2L0abKTGR7HHr7PI/0TDYZRCYhUsww1P7sOsMHWtNjG6qBNr/pDDCyaU
51YG7xiU5yY11EV0RtgpljtKIzgMTMq9bkQdv4kMX9bPiYIKyDtczAOytIfrJC60CRAhFmpeuT4B
tP9StjyPgfzcDChzpZZKu7uF2qHasBNKkyFtJkfx3mxxbmdZUkFSCsYZVKeIyLn9BMAb9WWGUesQ
3FVE5Ay8pT1BQ+LafkG+g6ajCS/81VVFovc1Lh7fTgTR9fHEyPIvT3xLQdUnZgnDr11MF+xofQk+
tnspYHZj3EbRkeNijXNeMDQV3qNlmiTOxguI4H4XuqvNNbKCMJI7cDxs25eqAY7aknvVNK6RuU7S
ncURbi0BzO1oKbQ9u7ZUEAUFGF7B4lw6ANd4O/+1Mx2DYmZ4H262DDdmZpW+vW0qDMtNWC0VeXYI
TIMR/iwh+8btqGTQZSMnAQSlX7TGCgPLrwdUzs8CUX1UMgxpUYYJ5gboOzhOgb5fuaIO6Mti0pfw
S9Zj+AYtnmXrIBAZly7ENv9AIvFN4+WQG5WlDr9PSEg8FfLwj/GBKhOpW/TOLGbuj0UkrytERKVB
Iz6xESbXryDm3Rl4C7z8VwybtU0lW68HJbgpu8clApozykNYV2PBazV47kuxROim8h/s7Dughh8z
V02FTNNw5T6JDut7AGqWAzK7+lvxK0Jc/R/olJpBQR3do+0JkL+BRSIRcMq9MPGtPBwyOTaJvXt2
v12JLRDDvpDgHO8bXlzdWfl7Kk8zsx6jjwhKs8oDyZTLBHx6EV8yp8SbHs8OkgwCLfHjY+njSXLL
V5G9yzUpvCAG9I2yiOKXmufZbHeObyiW7umGgCvW63z0UuPZiSF0vlco1nTjuP0hjlciR9NqFqOi
LKomjp2+C+RllRHja8u1DvGVGLuNPBwMynZjCspBZ4XfwUCBLQkWMW2PcJsr360XrO4J4QR1tHMW
QK1pc7c0xzpG4WWaGuXNv795xD9HVQDzOV+v801awe/vvD62/juarf06TVAbUfcidTi2QJh7BR/A
IwFTBWy462o8oc/vSSS3bqFSNhsO2xgWsambwwjxpEa+Vnq+0VeYmv3vlFpBb3oO3JI3T1+HBipX
YYbvjpNhhnPzTqp+uyl9JAfi39BViL89ie9UNlC4ON4ttqL3a6iIg4RTT6rXCHId+1Ucu7X2CxLp
79a9fqET1hSFGtqdGOVREfSVGsvtJ/1PjSG37nGc1e41TJWg683L5QnDVaYxx/ueJtzrSq22bA7N
MvL83eoo4fGrza+jCd8Ml37kgL5vTNHPGrd5MTV829AWr3cZjmC9PtBG8dDY2eH1bkAdY2qZWz2F
oWbg/qKdel5A7T0AXqaIkcfumA9mXIixmFo1+sm7S5siodZ1YR6v2KH16gXKSknvh78xb5EoWZys
5IRZPTKv99SHoKw8nkQ39WBdLKWqtsp7qdvKVxYRGhpUKX2SN1t1GF9LOf27iMzqFOS5p46ssIhb
4Jn7A+FRbho2s2ojF1gW0iLihggB9M4lHW/ecw+C8O0+2onhW3C0hu0YCj3T54hvyhIdb4Wofv3L
FdS7T7YYXmY0Q7YFnnMBZwzkI9dfJ3OGY2/LSwWLQOp6W/6ED6Vz9BoHB/acnSmbfx/ag/Ycv5T5
yeNruppUi2/F5Q+npXNJCg+3YGerytLMYAeaL58yUpj4yrQlOlQGk63GboTDQPks36+RldEqzZCb
1zFMn19W43FAJstCq3Opsuqy4gBGp/TIOXUo9xQ2qYl+0GMEaohcE6v+1u9bWDrMFmtUOcn9R+47
MP7g8CE7uyJSeiQSaSeiLBf4/TUzfF6L3h4xGzMDSRzZyfgvECCox7X5n13ktqkLd3BDYQehuTIw
+nvmwKmKCnS5FWyE0uRGbQwgN2tWan3n30iEUdGcRpKNMk0V0CenMVRLVhQm2gXawtKXItJGULGT
jDqW/0EUiyWkFKUb+6Gohtp9P9t4dYRuNnGGyAz6fdM1m/7nCUcFaFSZ+JwOSxXxAPqP4vDt6iOh
FTQMKSf6XP/pC8aSIlf/LMdylGR6h51qjSbiRhrGmXkiCa/x5PwhcsV6tsskej3Pzuc4/BbOakA3
18WwkJTaAStJIKYx4Mdhp1JnuPy007M/4nRGxu31aFgqtY4ZU45crLAsXy5Wotk4sbCzMUkMTXJC
M/KO1NSCMyPNF0u00gLo6mQUxbzJjUHTelwLYb3nOKm84DFy1z//dOTqAWED88/uBmScJ9PU2Krt
ZcUqbtN70qTyxyysu4h6j2XwDiylesjQVTE0VhJ8oQ+J4ZAQ4VvLoC7EmW87h+bbmd/4pvJVhIyq
CkdrjPuyVGWumWihZsQ56Hg1PIA0N2XZ45EqO3H+oJmY/+a4oRmznz1g1UQLMWlH+tagFI0Lvoww
goxcBtEw2Sckt606S9wowiuKqEGl7AJTCAQlZyexJ+jW4zyFnztOd/1B/XItlXh1Ulr9fqxP27i5
XEvTL9Q1RKz/4DgKoY8tjmK1R1JXX/gi1yV11xpremsb7XnaAac6vyzDXg93wkAkhA6fPv8o3ygj
KFtrNTazP6IIl6b9xJi9n2xt2wRzY6vJhffAKvVmE6sy6k3WeVwJ1+hBsQgZtgf+9xI/60xBA5+8
vxgtbpq41yydDSGEJy1IEjOAYgBOB0etDxpsErMPyFAMJB4Z0Py9HIdN5pwI7MVINlTgedOtrPPp
eoMbx8EBDz+VUYBASauQgiWm+9bA2XGgwbrqGpz9gXk3ZKeHkf1X1ZAFT2V+lzRavSJH97yaCGJB
IJSgUJci1pJnkatlSDpt2/c0PKU4yfqY3/g5bG7qf3adCd4n+yW6QjCXMtTBTslHid4yMWtu8gle
BlGzFuo0plyenw1gYdUNcD9/yTOfJ99y5bWXZCtmUj3Ry1uBdCa3D7WH/VvKc5GNOZN+vVHm3kco
HnzJWVX5x4knED4/2lv4v2qH3MIvWLYmjfDgVXUm05ZacctA4GzXcHPYssSaVAMcN1P+vy3biZ5K
n1MBES1EQHVlodvGZEk0nwYVlz4GypRNKeStNqqY6X0EbZGX3sZ3NLsXwJMrbZFwRfqk5QL7pqFN
2wrLuJ/UJRv5TQTY72Dp2wmQs0NGsv6W7zwIITe4bTH2J4RXjkIb7C8ZTbS/iJpLbmuUyvw7QLjt
aV/asF0EBkOlDKlpxaZFM++Ch1JuSHawYF4ribVL4UznlTW2jWCtZwVwgfu6pg5Jjb2uXn3GsH1y
oKz8NJNEgMlF9FnC16QhiGw83t0YxbjRF46V1BtiMcqaeuH6XOrOgug1qfm3I+Vg0L+ctEZXhpTD
OUB5S14W6kenjsCywJOdksTWskf/ifa3CQhuUbjPXKEks/d1dXhuHEDGzDPteLxtAJCwxzM35AOV
HOPmJ6j7EYORPJyPt4DeccKt5HlIX1NHyQJPDws9P2HAZC4O9iuvX1J4C5BPR5bmywOUhtal9Yrd
1Ql1t4YGXKWOTECJRPHiw2zElfwW2ydoDdDeLCUJXUY9vZZJ0bqM8LwVgWl1qoqaSmOV0hYdtlla
XXIDKd8LArNAmsU78TLFkBDfURJy1pI9ed8GQ8mt+gp9imu+o7RQNzTwoHzGAtbSPhy0INBJarEW
BMpDH9fAQO8Ltep4qCQHrIsI54WiLTh4XYpvOcMywiUxCLOlz5J1efJ3JaOA/HiVS4NwyD9JZ5Zs
BezClxI3RdnaFpwOCLI5s2uaLdDLkekO+53OkG5J8xtOCniRmcbq3RK3Bd2CJEKO8K9f/hfHRQkK
6jtNhEmguEXodVg0Y08dYyH8ZbMyuSsd/PJkax9tXgGlXSwSEpv+xxO/4BAiTiH1+DilPE5nUI89
RRI7cfSD3vkHTMzcg9ptP9EfPukgph9TXGJUVvoL/t+PZJV+F0ttrJ+uwcWPlUc/v0kuEqsPUCeS
ZJG9TqrvILaOl2oUE538Jcjpw1HjNSJAa6yfWTQdN/Z5Cq4T6tC6tIMqIlR8gZWodi4EPmyRNmg8
E3633N9hLQfo+OSysA5+lZMOGHFPcQ3IaFSTBKs0v7wUXyP+yDkxPFls+rrx0+cQHjkfUue1GQlL
408GRnhkQjube/eIyDWxRPr+XEK5YtiVuvZKKQbVRDx/u2Z4ZktEbW7CKW/OIs5A1UjCT67bUJkT
HCV1G3KzqU1Jbh4jy41nzvfFWWnlWlN5rTDObLIGgT3UoommNX2FsDaCG95CGjjMSYPUqr3u9HuD
x+oTkf2Je03SoNQjHjH7CGe5SQ+EaA7d5SRzE+1DsHTlR6hVAtluoqdbrWDYEydqI7txycOkenmQ
MjN5LzlHWHtWpwQKZjM+CxaDK2wnL5VoItQfT+xSefCAR73SHK+XlEsWvBn8vu83dNJRiBHFvhtG
OPX8zNRrv8GV8dBM+/+QRVD1Qh2xXTGsvYIDo/Sitr9ZVyFet7mY23kppwQ4KGsWkoOlF7JYgd4z
4wCL8zbwxSTLdhUmuS84alUZoTad2LDhulyInCQqgRWeHNnudTIGdGvHVCqTzRNtmZcc4XKXzygA
triI5aktT/qEkBah0TlSNiiuA33wsDF/igMBc648S2KKAEKcalDSdV+l+EuBeYLfkgla3pSTzgv1
YRFfH7LXvgSuaR+1Bf1Fwx1GSyDvOwuEa1aKeK5e7BTtRfiVoHH368SqFvVxoNkZbTY5bKJDKbZU
u6W4WGoFL3KTLzYOLQPs9lWD88zO9/XhupVsMn9Q53mbGVrcEKrRXg7UX/lZpcS9fiIdqkL/wbK9
6sbFK/6yPZDAuupcyB1DrpaRcb6NW2rvfv7ID2jqu4EEgYT2ovY29JK1c5EjstjBqxtR7sp7pAGP
NGEDcoR/i/SwpQaGc5qbB3EmIArpK7BaoThtbh5dKeclRoa0YDb9Xn2qJ2sPFYh83OLq81xVzQzM
hLXT7kug365I0Ok57N7FNiLWP+t+pCG9/pN1uI07RDPE77UOUbLaUdMSZZLjbJFtWHWutD3Cilhi
KmV5sL47Lt9xKIE65vQCC3M7PGNsTKdG2vt8lUOfhpxqQx6khvObgAN9aon4wdYVjBz5zg+z53+r
B9rD3gDv1s+w/+zqrZ6xBqkKlW+/qt3AVTp3pdIEctOrL/u9ier7pXz+g236xbfCl32VSnbp0xee
vRhSA5TimnjXplIVd7o4ZL1fzZEJ9ncuodiytBroJTshrAd6yHSSqc8/fCGQgdwKL+w2e5btkqQz
2E6Az9amM+nbcbWhd2s58RD02qa9J2D7A8jnAFjuWL/TrchtMOksI7p1mTC92ib73+ZlKs9AYz+4
jLsP9PfSpjgHpDwW9EPF8t3l7dBI95XWi+sMJ1A5WW61Kk8Yjbe35iLK4GAUPnTkP+k0i7IaYogb
+nhE8aPFLgaawgP0jDQLGw9/uA+bTWCYDp/whE4XMwGV7ju6Kumukm2YUNZ7yT660Q1pzG2zEZ3m
AZb78OnwTYWLOJWsPh4p2bWh+pt69s/5LDxFfjAH7FkvNyx61QEbaIeDjGJvd+N5F7puX719RmAg
iZ8g4pRNGEND6MFGWXg1/AJpj30u2lrJJcXR/EC7SUbaFouuOWsm0/pzb0gurWqvrEKuyAeQJIra
syonqOwsG9JGpXLwH/qo62Ro2zgJJIlA/7Yf5zK1AELfP/2OU8DAIQzMyw1bQjhb1qXqj6nyOHxc
abWp8olnCJlqq3yybuEw6lZylPJxDXpOhHynqZALNMDm89mWbRCtjvSBMawVEldBIPDjTSBe4DNP
oDW20dZws4PnaJRR3NPrmrkPdvYWzHcoEhsh49S38gjosTw4i3jcF6SuOO+ROl7Lhaq+yZli7f8X
3VR6j6ae+MUOPwUuuGBF++lTy3CvMq622KmdhQq/EwnJnFUQRa5l0K42iTnLvXdhY124nJwKmhdF
mzjQqtZus9kkuwS52GY1nnbJdKnqi3106ahsM1rdULeur0q1rfGFfLUtj+xpzySCkoZTTJUAT13w
F7MAymQ4alAdSI8kYJ0hnOY3b2/3YR8Cn5opm0cl/hbeDsA8jOywLR04xGur98xiNDx6i7Tod98j
3q4SX2VFCmouJjo7SiCRV6MXKdbdklsV5ZxLQaR2dJenYEY+jto2YOQh0ONx5XdJEnutI3yhFuae
QjEz0EV+sXCfW0t9a125jld/aGdnLXArkZJMZy/UIbt2jHy7Q9+q451I8GKM3YrBow4h15h26wKZ
VjDdZ8w78ox6tE8JCE4kP17rOexhqijIO0eW5mKA43EEct4XZZNiCG098nlDIyOZkdoB7BVg2DGq
RRVeQ/fCYwddvHuiTFKRiWIWsuVt6PSmmUJKcKk9h8kib1Z3RX168Kr3OzzM3qXBLA6ZZtpgHKZH
5CR33xcVs2lqx9kqKzHhQMcMJDsIGCw8ng/KHXdMMrMVlBJavgrSNvYP8vEfVCQrI9dvliZuuclN
e2O9bMUc0DbeDutFd1Ai+x0O8ZAKxCStPCp/4Rb+cJxKA9xQceQaEGxG2RJqQ8L8el1UtZcBY12n
H/REqDPelP7otm/V7JaGq5g6eF5Nz3skPrWqHtb2CDYiNnIk4Z/O928IcA6fbIpHtLxUvWHrWn1u
jGuVIfC01su3FIausqMR22ftJSKTe54qET2f9hStYARMDWK3Fq3gj6R6a4NGeVvNfjaESexbiYPX
Bblw5TaxKq39yyPLOzPDpXeg7Ej+V9QJzBZEUe6dyLvwY22Kil67iB7GVk3mKVcbsmrGx8CYFbza
NgviTgk0IfTBS4TYAfwU/nP/6UgH1zb5T3bbQBHuGHuSgRaWoPmDMI6h39v3FvTrAj55vJ5ldykr
bd/aXT7nU0XYG3v7Exx0eIcu/6k1S9UOUEdRw9+Vd2fh2cl9udiAiwOvKgQqVM/3Y4XV3KaIzJxR
0EOzXPW19Fk//wpNS07UPy2W1fBO7m4mHIHiytdzu5U/VUmlxJexRWb7+xD0gXyOg/9An0KpO2Dj
QhleXPSMozsPC4GXvBKGviYD6he9BZ23neLXzQW5rGNXch9+G8dB3o9XqThqn1UhA948H7XJYpAT
K7VvhJif0819TezH4flH0CgKuPbUKxltPd4LRrax5Mm4tymH8MTZoqAeAxfl3wkItZBt1QLdHcsy
LAPK0O6YPOcUHsoW8CP/68pohkO2OEkGtWpS3SFbwnl7Nhj8MK7VxvKQaoIuesNV9aQ/1GOiDfCS
tnPtzh9xZEnqY07O7r7oSgDwtgTQj1bVHP4Dwmw8KkRtwlxabq/blQ9SOiliWmrJvyhWmxaH3kLd
Gz8nGIndxsruKPEDBjvB3t7E7T2PXQYhl6ToCLwfSXjD+wuHAtqJgICFD3TuufF8975/rwTISCrq
NZap+12bfxqq3csj7GQ6pticrv+dc8M8cOFzH+s3friry6qoSlpNRVkJscK25qPh1Z8eCLj3FAjy
IqrS9QS8QsNYQmsu8RUi6qYGqAz0N+pevakmFJlQ+d83NW3wCdo6NfNC7Fm7iN3+aTP/aB2UJfx1
T4RtIbcClOaX84Le+TkcIWTbMOthQ5jTmiupwiL/kZVOsA80DFrllOMKlhj24qM73sEP1YHp68no
Gz/vVM0O1qLBBtR4HuYv8+HwIKGzAupRrWbCCNeyjXNHuzp4S7OHPi52LyjGcQp71p1lA1li8zqP
OwZvaSk19H03/CQO5yyfMI4+LlRXRbL+B1bSRAUO6Ifc8jAL+fmsN+UT1IbJMrw5oej02nrBu5nv
5BUEApkDyBjoRWuIt9qRlVY1HpXC7hA+QMFfzfywuCTs+/+DMvMBXUTFiueWbDzC5aA1PCbGefah
rFpKHak2+7RUKe1nVovR1qheFHgAQVOc+GMC2ma1fxcP8WOHLrr9THEyiWGsIspDZ9UhbI7xb6Us
pZYBz8bSrOr80HFoGKOzY3/DbG8HiUmq48ZgPE0EsHdjfJw7hb+ADzPTddyrdkZmiQDkoIM5EjKF
NTldju4Wn9ifTTznGInnjTeyr70vEV8jMxvcUW6uvESJVyByOyg+2xwDBX/sOEj5vJrVi3pKKziJ
onV1bMoh/i1NQIylDS1W1dNCj2Sdq22CpBmSG+Y4MJAPICLOTmo3Vu9LppTGNjSyNoMvSq0XFWqx
Q2fjImI/m5rbWd78mEo5JlM3fRC1uEEQmARfOu/466gyczl9UE3gQkmKPfB4jdthi5ZTt3f5i8AP
PxD6w5Gs/3WQk0uPUlhlV58EfjjU+obvsRlA4wwjx8OHwwlsGi25wrj58OtzkWbR0BHzY/jVn8qB
mIa09cC5bbP2GO3xAACdKTfxo+QLNs6mwnsQLrbZDZXLk1EGgQwdtqDYz9+Nic37SCDDBy3cRFv4
B+FyAkyOC8/sQQ78DXBVBlM6yq/uxA4aKAM1ckq0Cd59YtMwY+hhNL62lrOAyFEA6vImEgfkvrZp
xdicKPYuaoYyau9iIxkcnWHJ0ZGjc3hGMjVH6oYOv9Qlo69i0l7PRD741Ku8EPj0U8/HnID7Lbyk
4z8rQR9cylXln7DG9NZcdku9gF6uHL4urLNsuD68xStPwXTsJKn2UhK4j7wR+vTNP0+xw0kte6Fl
tobFhiA7eDIcun4jFxGWTq0sZ7IrM8JaAhCuWo0Zi0F9zyCfh/N0VpkfJ7PmtvqXG5WlmTsXYx//
qaZT45OQsegqokLOnMfr8hnZRszc2fMd4iqRt2r+4/hXGpmUuipNXcr0yN4tcbLL3ikza9NILqCQ
Q8IMzJKJkUgjbzU4aDPGvONmXI/RVQULXegIBAYTCrmona/CidkZRS5JILzt1HPUIMz9463IfQUb
/Uj9El7dvzaJSs6+GK/r/9FrzJw1nBtqE4SRMbOBfcNdY9XjMAgGSZHs2VCkiXbFg75f3sr9DYrw
h/jpIwu71a1wPNdFEGK4K9lu/Jw0ms/NRj/aahjP68vvR16rOIzrohJ7Q1mHIOIAzNFHG67uN7xu
h59+3TrsO48f+x7y94xXHoWTg94nKcxnqgxAxwtM201E+oshw+cb6QCOdoudDD2wCRHN7F3NXGAG
iF5Wz9Cej15ZmctSLzMGeQfD/8HdCG4uJYO1HsKy/g8lM1waSAVwi3liNuywsKKca2rvz/N2dKdc
VATG7icGS3KpPRlUhyfYy02Yo/y+pZYq3fmvg7TgdW6KdSVQbXJGJ18aufGfOrE1x0VI4UtdL4C2
33wrZBVo63j7Z6i02vy6cwZx3e4I/zhkYTPznAZJJ0jnfr9Wz5P0GAIkIkAK6pH70M1jsj9u0JyG
NacFAKx7uYc8LUtfcsb//WljRnHwp6ul+tiq2fZ2LDQ0Q8fG3W/jvylTEU4ewHYx3mcEv+sDllSy
mNDWzQrQzL4k/AhFAM2dECU81hoS3kS7B3ykCzhnDpzgR48S67v7xtkTLc7drF3MNFP+qjg6l2xF
YKD1h2I1bFun00KLOpo1eCEpsNTbsVIX5Jdi+7uQUopUvaEKgB/WJvQQsijspod6NScaAaD0sRa0
5Ewk57I6BYGN8SQbMxTvRBtiAkydmJKEWMZyt9YzRQhKko69P9to7m4FD5WqwOwt1snlR/1eJlU5
tcERWrQ3aWBTpX3hDBWn5iuQNozOt1bsfRZO4ei/CdbhlYTJ8MpcXSyBwZTDN08siSVYtLuSan27
PtqDn+R6xfa3BpSAl3OtTKXocchsb6ms4Tjc7RsksKmNIZXqxJxo4kuVjSzPI+X2MgK6Kl74zS0l
EUV7Ha3LeaN6jrtchMpFdfW1NVysyw/5cB2ikwP/589yw1DCXeBuUCr26qv+EYlKmz4QYIXmHjb0
LpnsTJ58JoHDZ4KzlpgMl4vHHyRaeaUSLkMIP+QIBifLsSxEuQvNV9aQA6SV/kRaMU+OZG7CGqRl
5GyOfWRH1A48M8IAQLVbkX6wgjexquHFfa+Vaj0pDixM5DROJv79yxPfpe2L5bwWaE2Yizmayt7L
nk5wOrmqti6CJKoIya6mKSlkNKkz4JHCGc/FClNbG7j4eJY6HU0XUeSbfKcydUPbqCcqNIKghzaO
s8yTzDaKcJUvJnVvd+2wx0YImDaqo2U24DDE1jUDKodvsBCdHHJm3+SWqIeOSvDIYK2LEyJqsNWE
E+Y6Dexr7AUX10Yz2qvKCyJqcbmF8bqJO9PaD3C94daRA1lOL7qJjd0bn5qTL7sLubxJfD0AieLD
scW13gjNMFbxcn02cMFnpK+o1Ey9VhAcDDxLcXVkcTZjXj2ZYPZxv53YTK+sWWiYnSynJdJ3ICje
rNLHCoFpjAGvTeHqm59nRL8M9cFADV8U0FZ65kuqzLcBpb1wlmK8I1cn9jh0PJOEROPhws/WJJNp
4k/CxhG8cM0jnXMoEafZ5qE+HO3afEEdtVWK6U8bGoFwQOODm7xbRUu/i1ETaLCw/0NRQ5syCdsc
1qPNXale4562k+dToHxV/MEMOaAw1enSbrNhFyuEX750sDot2t4UUAkKr4cMDk6K2NbPQTXjMHs2
hHnrPeSlV/+JYmAd7xVpXVEPZVCzZE2lzigxo1RSiwyVi7DQHbNSZlV3bjHbY2g5adB6ytT4naKQ
+ei514OWv5zKnmgCMegLe8hXfe9hTwWY++6G/dOl0YkTq8r+5oNZCgxaNDiGRt+d2lsRwcIizxis
y1NS5mhcJPmk9vY0hRp2PfuJTWD07AMG8eauy1iUS5h+SJgmMncTGaxaghZpzDfoHI4KRhG7dLDW
jrXVqqJTZlmxrwL6mPTBXeJR7EfYvBp2OzyzjUvt54dvOZ96yI/m3QRzHoqFZVIAeupioERogRCT
XRnGh17ZnKgIBYHzWheuSO2pQ3q4Vrryqi5IgX6rAs3q7iL1O7QyNBUNeJL35QUkhV54I144dR91
bvw1z3luzrn5j7+4vccf5HXsecyYjvbdf55A8Duni9gxpLO5JtUb6xsHMF62p576PD/bY+kUyV/l
GepYSbJwaLXHaswCK1Yx9Xm2TTjmg0G/ttlrefOwod1TeGk2bWq5ghy8Pia9oNbORp9nxTLb4sG8
0SW9WvVAFuQhySWXGkABo8R55Htl+p+YwGY4/5wO42kIxHzyyD0qcEdc0Uss6w4st0Kk09aYCLyP
cXz2+WJQGtfrm8g/OsdmaVkt/flP8DTNtTYk5PY+h2ns5VDfdVPE7CsrfYc39pn9OkXdrKG2F3PY
4k9/Nmyk1JyAPmjVbIZFqan8li+pIpdtMhea15fTT60XNxtyzdNxCususAf3impWQV2PJdpRdZgn
kR4ODdl/0EuoEtPc3f3AGfpvmy1v7hsJI8xZJpgt30yscKTFyimmvET2656/Dw1OE81SbTCfbWOl
ApkBzHlyC+1Qz85oqtjtk5VMTPl6+2k11y0UO94uaYZu0Vl7qiB1y8EM/zHKkxLPQFFFSU/rKYD5
Zlp16sSz2wkaARJ+Zv5LcLGmVr6s/jd3mRT0Uxd4auCBb4cPAN9X6vd/2m9W5iR8XtX6pHSsfKDl
TDRMSBLY4e2Pcd0mfiH88ACaoSBBXHYhUwLeJI5dqEohzIhjS+jmAymvv8MoCxByaXE8BbLy5WUV
3u4Zdh0FwmgrH20xw8Bwh/yiV5ED5Vb/ydukdy6N3DU0MlYDNR+KSDwAsKXvRBf0grOu7Bux4pnm
Tn9Sd1h5E87Nni2WNUbiU5fTIDhceK1cjqxqqMnVyRi6dce8xa3bKfzsCN8UlAzLKFbTtzMwhxYq
QS3nx7RHkashEZGCnxcB+vA9U9iP9CjzFze8sIHvYsubiD9AMbBjfdqOw3z/UkDQ3lcMFgfYMm8S
ZL/R75llJeqD3Lvx/epyfLV/PbdGxjgOZzQFnpubtjL54FFTCm6xNKgt/P9rqF/T45FmEpu61Y3L
w27VZ65V5fY+Cf7fRizPJ2Ab5+rEbZ2iOaxPnzqx8T+1wE/TgRSEuugehnTMVGKo4Za9vJQ8X8hi
DQ4PelaR4BdZAABQiCxd16HM6aYq8XX3CX9uGNLM3WQoCdCVxBDPKg8vrFETMe8lVWzYq/FQIAoF
tlvCsnQ4L3jWpO6L5OokXCiqPf7OcNxmusIG7eVtC6gz8KI2hQiF4STowdYMlSS7/GYg30O84Xod
ZtjL+5M3CKYB/NTuBMdDXnrTlRVm6DVZLk2euCgA1YXbjN4fR14LS/YEMHuXgV2yr70APU5gbHE+
7W01DG3VAO0oPwrJS6uZ96UBPjP70a8cq8+8U7GY1aYod6qELKt7DQsPjUtNS7On9HovlpKnu0gQ
GiVaSPabX99bII1MR13Pb9crOJ2qhTwSWKB3sSN4t9RNugq1DWKJPry7zcbH0Urwvs3XRA6dn/B+
+fvq67vgh2YsWTMpYgBM0xLgckxZnlZXpshEsfNalaVXtUXQAVp6XyrHBRobCGcaKbSvjwU75uih
NBAW59nnnLqRp4PqrOTs680KLE+Ul97LeTD3o3oIoTOqLmj7HRlbTx/UOpP4aEiI21cKw7AH3ygn
BKtzsi4iEV0wNZ2nsQ8p1b69jeOvGi/1cRNZGIeGYYeYCb5JXVui2s5coyiBcvq+LPBvp7V6u/YD
wzIBxfBn23IP+RyO+SHO+9UBB6bHZ7cLML0x0Om4QTX2SnFaO7eQXJW7XkfuYQJhYEyD1jmAoRhV
Ny7DVwUZ1FJuHWeTof4nWARR70iY5nfTksG8Ep/9bVYzoYjjik3tzWBtHXzTP4AlNNfLwNhnVs/2
mSJNOjTOUX5W/UM6i8qSs4rCEezzoG/Z6PmL+wdax3o51jmzKPPLsB+oCshjSL6SYYOLsQ5OL4dN
ZHYNUZdhZtFjDc8DuGaHG+5pgKjt5+4YmJ54w0O+8kDYQdrqMMnOeI8JlVAA+PW7Cy+ibc1ROUNO
81Oi5n7KuL9vW87HMKI7Sou/gAcAlmRO0K6z698Q1VFnWbEWfGe43MNyK0x7HusaO2OoX8jAShEF
0M34Qv1cl9NnjBcBS7/Kx1t3EOQZfXAawE/VUexj5ziMNlrWB/DAcu8OJ+r1x9I60mXU8anMr4Jf
YO53IrK7He+b0vXx7PshyRQOI86BDqh0g6zCFdc0Yhl1T87fnqp0qxGkyj5En8oYlI1DBMVuFWzv
9q9m9uNceRn139jphRjdgIeybqqYvR/Abl/mr+FpNdjsjUQ1YauilU77ceBCRnHYxws+1OM/Jd/P
A4mbsDjMf+6V6tEFPwlUXvPnpsA/1IRZVAi70ZUzjWMG/9xJIhOFvt7/U0A2FicpgqdQL0Q3o7c4
E6drEubfM7lX2Rm+ettZfbqB5RCzHSdnwwYSCQOV8MvWYh02O2KMNjYi7ZoObkK1OrzhX5p5QjS/
aK2eT5HnVvBbKjC6OSfKVnb7ofCHQAeoek4Tu4+H5xVkCPrVXpvHAeyGrN/XhYgqmK8hp85vqUPS
xfMt9HIrYk4n27EGW5WhflxBPzbiRjriIsOuOCgjjTgk/G7cJGNvQRKFh7bQcDSJ1HuOUkOMaItz
22RFtEKdEckYPR1M/ZZqEjGygI4imX2oXhsRZDIaVAIwYWuaJRUdF48fAyuY+M+RKCt6Qh5Tiawa
dEax1GOQ+8o/yINMde7BOn0raWim5++r4E55oogf/iGRbZdTqohMSeiC9IL8CB/PcK9UOTMeqw8C
Yh63aim8oJh/kvT9KQTQvpGsItcVYi3B5o/rNVc2VgmGAdECOxnCuwQ5tq9gFOntbgPn6u8MZzzH
FWo0X4Tt7FAlJyMMekeP+P+1ViXubiyU5PDIJXSvuUrr9jHApT6m0GzutRXCt7VnNQHYzpU78rZT
aQPuWJfb1BxlzLNi69E73rUaNvNYIt70iYIVpM5KYKrQAjGYh7s3ivLqDqj/oke19NHvO65k//lA
vUHlPeENcZc8dfdupTvqNIvNUqgBjq2k5nyIb7e0V4kQmWLGI/tUlxN8fYFpz/AGyc/gnHOVhU7p
dOKeyRyDf3V7GKVkCxmIK7kfRGPkrh3XJ01japTlTgo+wd7+sblY/ybo2bhO1M16gLHhLJNmPshg
oD8Xn1iu/45eeEMMQ7DPQzncTAe8MBJGMrcpokTmmDk0itxgW3NhzlRvTaIGxjpsviBJciESRqOi
PZ3cWTkJesu8Xa1w/mWomtXFSVq0SemEVhojUT7K1TMF4C0bIgomOYHaBRMFBzGOX/zkFDn62Mv3
7IyWM1PGvQp4md6SQimHyIzoscU94CySvaNVQqksCBBjcna/hsSuA9ldBSUASpZQfRFgnEfpw2UJ
GvGAiViRMmtr+Nv9AyTHq0N7FSiIpcUfusipS08HLEcNggqyZNm4e4Hi/2K/P/zVuJRpvOllGXvw
2qvzazWbG6LOE23xQbYAk0++O0Hh4hVbjYX/F4Si1CIbvLL+NDrpokInL44Gn5hYfU5fU8/Rze61
4kjeW3oFlkfXOSTFHu2CpzVNq+E+OS5Thc6W7Un7Sbl7JhENqDmZ15vz7dHpWK4cG43VaeF4Cpn3
InpVHgMT2F2o4rGDUHh1fkz+efjF3h29N8MaPONW7wXsic9L+xF8OJ5SyrDpg9RJO4YW04XM3Ea4
Kl4pd/Pl6GHCTSNTX1qlkQZ1Do8ceXYgRmSFh4+ejTZUAfUTe1I7pxOqe8cPdQHfKt7Vt0Oyqnog
uTWTOHyThud42RDzrH1t0ctzqSMIz9FgskPHLdilIS3GXjMLb4B4WJmdcs/6J0duzP5BbRyWr0Nh
Jv+kO/a8+UNBSErQv3PCsJoNQHNAy4Be3l0U/+KhgTyGB2SsJGSrLO8Fk2vlJpU6yLGES4IEPwPI
jPhyRNrOtaWwZL/uLEMQQJnkPnDic5SBcHpQoG7BK6q48vIU7iXO3DQdQsLx0csJ8wrQOstrGSvd
uBL3gc/VPXbKcoFIMTrPey9EdNG+obSdFDUqeNH7ibUmZD4E2zIt/GTcbEqnFzdE2nV4IN9zjQv1
2umDTcEOy1gRBkZNMxp9PW+HEV9BUjNTRAXYC7fkgTl6pSTBNLQic3nctq3/R3GLiQK3YoUNbP7g
G9wfRzo6/npxuQ5J78goxyy6leZBORzAjxl5zW1nOFAUqxSunPQgWHfTTAENPoi+rrIizMROjpTk
8FIW1xsU3HwqQWWt9blV1nDsGT4jMYN9uxvSRqHkdoN17IqIGuMcClpI0yMtSY/yW+zTG8/endIc
chg1fkpTIyV29Bado7Jl4LlaUgbeUHePJ00sBUp/6qkxqKPTznUyIIpX/mnqXQf7/l4bT6lb8mxh
9mwrDYFGZbJOSd9ZwBDqWdNoPKPc7cV6FshSMKS4ABHWlRo70JK9UlZ19uqzDi15Pph8pBiv9WsT
zy7OCnj2ugFsWGzBJ4SklvfhyzkRY/TOPJtSDwXYnl1NX/+F9n2jRJsCQ60cFNPZkUUMdySAvhxJ
QrZk3l5E71gN2DPlN/Gkw8bmL5FbJ+y/gRC23VpWs2Q/N1OUodKCrMsugfghwXDmgYvCod23cctr
RUoSnWlZvvUCeaypFEm67Ee2KhujRO0bYcKP0BhKAAMIbwyokI0R60zUjDs9wpsDjU9AsqJAUbdp
Pu+dik6vbDbIAbPx6fHIiDG65A+F+kJKBhYSWlRq79ESRCFNrtapdp7+GITMF091VEuw/N+6AjDo
GXxF1XefQinlbCqCRLhYs7jyeNLMxHwL2+VeKyavenbIGrkTyjr+Zu3ZnV4axS0t+ngGznPmOZWR
beCjUOem4OcVMbU3uz4Rv+eO2ysRTS8wP5MMffcXjeLqv3y0udIIsOpE6qkSfScPuPWUaJ+/RoCt
2V2LXsV4SB9nemI1vzIl/zthOwKdN9LpyLowwUUrnK4rrX8pHqD1n0i+sdECjuEVBFisLJ19zH2s
qI+9FQ18ZxDB08tLVEAoUyn/OyyoxUI+6uA3wA40kenHM/i/A98m3yn+IYRd6ptXG4vyeRD8r/dN
nq1KlM+HMldz2idAbSxMmj7gDw1VOlwOi90jpbNnnTEbqtQ/7MaCqqtmNFjp6fCqxjo0SpFVEQTJ
yHUYc96jwuZYUvRH2QFv5cUvvq8FvMdtVuthHIAA5IFNVZKmw+wq6FpKPoI5bgNjGskM3kkI9eh3
IynXOHbM9VkdBI/btKTsOxhMJHXj4UtWHYUv2s6oSXp3YX7KfQiLCGDKhxZytSDzFOyFv7X/p31D
cDJg7JT81KQQhJ93yRxWFq7sQFygFfcUK2DjLvnXCSJ6nGr9EUoXO5vmT33WaEyQWXm9jEKtfqkj
E+Tcr9ZyPb1XnG287jJOrTI194lFutbLyaEe7tQOw7Ry59ZfDBLJMW9zvX7+WI/jtHtXnFecFjK/
Y91opy6GM/uLrU9YI8BrQaZuVyBbHgVkOcE3VPD4ggwcBuAVwaLIgr3OxWDzKDcTrBph60BUN+uL
9Dw1mP1VMxaLiHqZPX42vHVg59QsuXlsySYd2Hn6+v2UqV0l5ACLiMk/3X6O6VgrpmYIJv37NEXc
bbazFlpPrZeLvxgvwt5xz+9d3dP1kT1OYRHrrprd807t5F4/WLm0wY/mcqNy2OoT9zO1uJY8NZAI
a+FFheyRgsa19231zbiNuj+WQn7W0As9UiE9qsbSsZlcQJUzswkchsbtdu024e7C4sQYG52mIoxF
6eN8pxkBdrTz1SFdP7iYfb63GT1CI16ascViHq/v1q5Da1yMaJXILlllxLcWL6sm2qQs13Cf1n0y
Kkwpmko3VQEWGxykOHAPGQd7nJs9vC9A8lFozUYLE2Kqx8z7HsgWlfYa00uKtPJUjtBnM/YRea5T
rrvWkNHGQz63DN35w6Zj6MGMtkQiSI9jPH1v4I9M6od4X+FJse0/UzRuaYzH4sUZp14LLlJJ4PX/
xYFnyQnEs7o89gutyiG4adMZdjC15wXN7DpkCDFlTSRMabxA7Ex2j6Im2VOzjnqRXSS1QbBqxrws
+IdfxhJv58E9AEhOMqrNNL8zuny/eKdV5b/fr6MLMOu+dOJOoyn35v3MZp/RPew79sfb3GikqSEQ
RhGu24w/GNqda+pCv/h+QKTMoUrJITz0BUCA10vNeJ5IDGvjSHTLEjqlZxHyEUnadmpw7pfaTinf
nMxv/7cl5tvNbwrFgCet4lfn2ze3qD0NCxL4VFacNsJi4N/sX3bnk+mtZR9pUJq31gbPGk8B6qth
xvIVbwCVhTPy9qKbKAa/9LCLgNjtr7MjCPZt5NvIQ3VF5x73h+UhgJXZNONHIXjp9XfPC558kC0d
U6gEBz7kITlhukAkBD4/uSskzNL6DtnIsknL37TqDdxb8uDF9o4qUDGgFfyOAl6NhHcRKDgq7e4A
lc7PhN7M7VmiHA81pT1Bgg01O1Oo7D/dmCa9G+W9Dz9CCzx7ruQurY5TcigwUCiR7RD2R2xhM569
gnOxuTOtuZIlDD4GFUA4eeJOKEjC25JmUmFGT8/AWtr+7FKcUcpPSV00fOnhftscu8yLOLnwZk59
QDgi/XGhJ/icx5oQn3Umb/gr2tvo2ZU+z2huNeut6FRncFESYeFg6fO8p36327sercYVVD76wVky
eGlbi/bXmG2kJQr7OrIvZ31ZM/qm70gzseF0Bu4xzDFeGZHJBQy+t/xqQUDgwk0VjkeeJxvD+2ry
3wQ0DMu7t7PizGFjB1gQ9BED9Mgvpu2L1aaL1wfn9u5N5uPR//4scxKN5z+hbHW+09ii1Nms8gAs
nsCANRiJjaBQILp9KPbR9zKe5o1QozuLDTTlMF8lTWKVpNsPCesu33fW//LjoLuLyn0UZNhnMpA4
M5RqQFBhJwddU1ooi6no9vjAtUTPmV6iLRdJDjiZjFTY6MV3qehnRwsocgX5HemhX8AHaJCxWK+r
BcjynGHmVhQbgZA/KjkFQlWlknQpXD3pj+1ifA2MieG6xWI2WZBbqiW9B5xRgAe18lCLlLPxgCNE
XHA3PG8VWb229IvB57UcNmu07TO6QDOjnrKoPAfXMc1jR+1rTa2qlGAfVHZdI28Zq7UOvfZV3we8
q6lb+7lQ1j42gbNxOoldzaWE974MQ21ut1QjWFgNEGo6q0BKVr/GH9cTs6uW3JBewLTR1FEyTebj
mTudraeIJflzhu9JpTYLCws/Yt+vp0hdt6SsoS80Njhw++1DAfYn4nEzPexS1KAxv5jubSon0jWK
PhTPzhEwtXtLMGphdku28rGw3XK2DUpqcf2ErGU6Bk69WF+eGbQZc7yKn2Hr8ZaYhkxX3fTh7rR9
oLuDC4ldIKzrMiWE6h+r2O64N6xCyE8ic6rttiC5x390s/ff4ibxyl9Y+qiLKonY3hUu87DyfaZj
er8Df/Ooh8d3CaEz3Sis2JJrSDis9jLePvXuzD5+JqbLF4kPkgE5hHQOS8P+E6pFkLN2B6pePpjr
KJakUGjI/KPmz+05gMVsLFmx5i4PlKJAQedJsGtdRTUpKHyX9eWUUNc1bvW8n8jmJuviXIvCpXOp
QA3lzxSecszzERA0vn7KcVhilEHII6c60Judq0gVlgldFGE8K5AcfMqRJ7Q/riBZPtS8uIudDyDm
wld/Th9arVlWRpuc1Y8RQGntJUy7uK6POatBZOfCOCagVFOXsnV0/8eVcmvxUI2h8PCfc3UjfHVP
ZOVw/Ayn68Spri0nrznFYTZkYktHZb5U6HJB9sbQrpnOQHtR+S9SpL3HOIVbgmY2MpPTs+Z+B3E+
EgrbLXR0EsxEuPgp5mqrzqdmxzv4SOrHEBrmAlqO56TvSbZAcd0Knc+Sx3JvJa7ZZSssqRihmZIP
T1D2zGKHT2x7q6oUz1qB4Vx/wn/Z9C5OFR3y1CEUj4M31McJ2cFESRys7s9vp90R6EWiChc8GkUI
4BJ8PHoEXFwoVqJr5+fJR2EEpgQm9FeOdGm20yS8BWK7o8KACauNgW3qJwmokhO2cHYUKT5zY4Nw
8cjya/W8bt3K7YhiSFUAAXVX1HqrzG7E1QlHRIJ6iREa822Wv6v3EWjx6FEIDUFSfetlke/3+lBh
9zCE/NfaFPJlqILnx7bmbbRdmWOUhMmp3gfb8kJ3qRw+JmUq/hmK13ptc4VZ7k1V8zowGZHJZn31
TutAI4J1eqQKxdIL60wl8yLqWMwVzMY5uBkP9i9KGEYcc/Cr9q7oHtOrY4vfnKpixb8/zY+MFSb9
yMrfB/87OodIL71u1Maq0OEzASEqQrhGslYz2xbUHWUIbjLS7AcWB/kaW0HIuFFl3EjfYQZDv21y
HKWmow8/xpXd9AnABo9u7NK5q3G1pr7XygM4NUDscFWUdnegKe4mbyCNHAWFTV9a2QoboClHA/sp
fLjz2Zi0ZLhaZh4cTEJ5PCUp00qEwe9mM9CrjPD53GSmmUObB4tf/Mgo60huW3JSrqtwe0e6Ffx6
TrkggcwRxXcWV94Er4Sk6vMdxVXS3w0jpyVZlFrZI7A/IoLh1plzTI9EkHgOJvyfgLy6Y0nfBDCX
DqZa28Zuzf1RM/6yVBMywHJdYDIT5i1kzBt5T4gH6aPZXDoco1EOVEcNa4TGAKpbg6mHMcAuNy/3
vMWaVoormg9HEhETt14TDYoxy40J3/KbYxj5BC1tFQK0XEPCx8RC/3fUWtLBr43NCwvUooSx2KF8
Jo/mpBOTXV5Y79xwH//fQPc7bbD4NC/K+/Ef+XMCqFMcDYC+lHyYxiW9n1u3CAkfqPPlPaFsqElV
YyppZgNmHGXqnreLASIuYMBPqhurb/SxddRBftyC8yWBY0WYJRo3r43IyWA6dUNmva+i9Lmu7fty
bjEcQgiHwHmm2lFGjKBkLUdTWQ8riItQW8EbXQ7ZJAlJIioeRqLHApmJf7jtBoHpBfVTL2eo4DSV
cbIBQbLBa2+vLGTYLm1DZRusWMoNhBzLrdryaN61qQYu+pjIrSKz7YBgTenSVB8g2coi59UpXfhS
0AP91e0wJJDZfQ4RC7/1XtP3HC37UgknWP94m6Bd1OYPXQKVKQuIbO6ZSKpq426sGAguQ8ZGlgsU
3n7rvlasPjir4n+NOFQAI0N40fF7IM/lDnuglx5a3aqjNDlqhv36GOXXYiRHMU7lTRGL2lPlHiNn
QtjO4p41lwANyGDtPab30+kIxKChaU4Un4SkrV8M7uepuHCuoaGEpM9LqmY3UGVJ1Ers9ELRa4OT
6HWuw/Lsxco6Ye13z2I8qGeF3GVOFjcxnnBfup9hnxWkBMlPiAjZdcEDyhYP+JhviPhstCUZU3TP
seWo3JFFjhGbGfp4J/q3AlX6/c5JmW7pOJvq7zrR7gZs8Zh+lqz9gYxHm79QuQCb1KQZEnXKbG16
LLctzboaOplgioit3Xb3kw6jgDbpjJdFrJIdQHicMLAUl+1um2p2MmzxY/Ank3ekGF4cDL4RYpFv
1W2BVsCF9keL82uXtpcXwtnMkXJsGX8pPfm5FGvN25EI8vraOrrk2ZYit7h2Tscift23cvjrB3aQ
jy9sP+a5zJN0CyD3bOZ+IJPQc8Ld3Fnjp2e5HYRfjDzOaxsJr8jU1CFWXcNz029bCiA3oqV4mvtz
2wQ4XUTXypkHTXt81xmmFgBQpcJQpNadwPQ9Dtp81Ux2uqCkloGLQ7yYnbnUTjwEVyRyZfFYxOAM
9wUM9aiAILk7Pa8T2JzG4ZvJ/HlBbX+G2TRNgQku7+bwcrUtEKn5toCQZ1H03ACilVz6ZgW/V3uK
g34qx+JQkt2ITvFLnMeiMnHmrYmDQNOAe2TYIrMvFpSMKNVXtBXBzNmZKOIVn7W6pZx6qIDGm+vU
rOB9PVvNT2gCAZGJa5uk5g2GNx6WkXHjMUUvWocW4F/XW9rk5nfyJii7lubdeFurg8nl5PViRFzz
yvv1iObyQBTdXnZO/zXbK6w0c1Il0L8/0ZDY2F1c3furU7ySyiEZBnuTnAAML/AEjFcR3qvYmvzE
HlEE/3Exqa27JajkJg25v7VowKdp1ii7n/mVeQvm2xY9ImMk0nF7IHWUWhzRxg2SkdE0dZIScyTI
bb1k0/fO9gREspIwj9AjXaWOr2AYltNchIAwIFMOjr01KpSP+yTlVab7vUO3Ca7J3i4I5dZrOgi9
eAuCq8M2l6NKAtYwIXaNACqLKcPsov9kS8fcJ7gSxrAEYNplYDQ44E68ZaWnPhPuWT8DtBWkVP8D
zYbZlR7p343n3y6WrYQLkUFaeRi0YNHQ10N2iqg2T4iVABbiHCbgSMZwEQGZ/6oI1PWLtTSVHPqr
Uq2dqDbsjkbc7gQN+s5PPjNsvnVfxeZfJHUTYZ+vTEmTNsMQ1Ldq+i4zFoHFKIOKLzesQ2trHeTn
s0qWATwomrsvYvoNnho+FhJiDuzz61ryEWrHY1rwTMHR4EorowSxQkuElrsK8YLQSZkpGvtmbG+1
xBh+Fr8t4xJArKKVRRdPrFUT8IYdW0A2iYyIOSCpK5XTE8+u2fukSw18nrKGhOCzWrqVrsMvrEbw
3oan9WDwJp98/1fIfJWA+X4YnkehPQ26efW1UMGdsh9n+y8Es8fpzANw+mB5E2COGE8+eowp7GHe
D8iXnDhuX7xQ3yoa/663o/26dtu7zppO4GoX5AsmKK3vW2A8Y8xBxFUAnn1FHTlmbKdwoGqQIB1S
ENiXBsdNZ4jmb6sNr5k0rtotzOzCSDEUYZTFKJBy/3eTzndDO71NnOFsxymdiRNnldU6dP9h2l+g
SkV70xyC0jfwfkvXmAKY765ttobIPGReb0hnSNA0s/B0kFPmkviHo1RPxSrVs0wWtD8byx15WJRM
+oXQhdGgaJkZw2T4QmbRInGQ3CfQ1HztW4FSmBsLoC0jJiiL3pZzmjgAAmDoN8PgGwhlVIViTVFL
ch6W6dM3DgDoCoGG5iUIB0q4TG8oX9gHbIt1vcVV7BlvufeYBJlhub6VEyqpiVd1NN169CG+90kh
TwpuUCuY66jTCZDdGCSxZ2ZiDPe1A9nWWjD9cYsXLiwEm4GwHPYH8r/kW0RyfFfikbf20xkAcFI5
bokjev3NjAMPo36pYIzbObku7bj00MEx7OHb5vAiYjqcXv+xlLEnhAdn3N6nrQlONfH7kiZUAs7/
9qLtepaR/bS0sUH6VP2eytcAw1CDo7pB2qwIc6ajGJ0X8yakKmvEkNa+KjzxRbEfuY4mYGbONJDf
lYnWu61Bh8qCOBT+ZRx4yVWMsDXZGJ+6akSaxeSyxXjzlHPBi6sDVcAgp+IJ2NA6+GLHVa3AcyV5
KdJNPhTz/aEynbP5gC700qA+90zganscfH9oNecbGkk425hSRzTT3crNKc3XUZ4YkbHMb8APoPC5
65OLNUYE4ybcxnXzJsMDiTdjZF+R8XO93gprOR7gvaMFA9wlJV9EG4UgLXxLv7oqDK8z2DLCvXLC
Z0v0IZlxUU/nnPZGxPE4fhbN/LPibOJqOKp5Fbpn3k+TMU0S7fHocZg1ivXbnFfCONzKB24vcuU8
iwWrsMrJwu4rjMP/bIWkar8VXrRQR1SBNaBBDvmXHShKO9jLtJLppnepmqh5VQ3Kxnd6hesG996+
uE3SqjTPYbOG4Cdj1opZl+RX7jhyrmO+LtlRmipl5mdBVwBy/SbI3vNjFwR0fmKrSE1tsOxU84Cm
AzzhqxVxyjVSKmomJCcCamk0Jcb4NPg01ME+zopfmhLRIaLJFwIdgWGN16HlLyGid1MD8XqeiE2a
LMopQAK/dnJZUB40GCqLXfYCj/OwsM3d65f6b6Rj/5VCzif6pKWXVRl7109B4w/aLlMaGHErMfAl
cH3p4Ty4A3fSH4lwBv1C4cDDfLcbcEkTN9RYPkZXUCsFUPh/DUjuTkNNN681h3tDzfMOmyp5uEHk
fDdadxu/cwyGZwt79u1MBU6sf7KOmdSF+vLe1gdrnItxAkwRnt2a/agAY4YrI4XZlPLhH4LuwC9t
UoEBtkHAEfEJX83wL9lqm1CwdH5NW80oiWh+Re7c4rTR1HLb8tN4/uYpA6SzLA2TDyURQXlIeAmi
htzQdN+8K/2ocLG/Nx2sJKcNBxvHwzEFPDGcVvPuPUVRtdPHLdHv6YWO3YmSn62GcWTT3uOZCPUu
NYJBmSQRGyjxI2w2iZv6Ich3tDHIXR+x0hsHDNnNMyxekTKK5mfhgxGsv1ToswrRxEmLc0XaVcAV
6wGe9Kc08dVX2OJ9DCu4HOyj5Wu3pzRmm6ssNYMqkOMP/1HKRugEYsAR6EmfvGKrv8dI4RyD6gsa
HKYTHo5Jy7+LdrNuRGy3OSlRPLqV0h2xOlNd3VcIpaqjZk6cQHTR1eBArLujY8B/y+6oBpPf//MH
OpJAXR4leyiyP02jgNvcP6nG+l3FP2GmpCdwNe63GN0OJJ+W0fhF2VJ/dspQjYk6GQxGuVEZ++zr
1lfq7bGiZKraEtEH9XOgLLt8QKS6ip2yMe1brK2uxRXdMciJ4apgdi32T7h7Z/WDXMn7auougWda
RzlQH6he/PmDuXT713B3pfm1tLGXYCl9iGKtsuPCiJYPK0E90EK7f2M09Rt4JEIqcYb833hchil9
cgin9kFVYXGvBFRiLol8dd4XEZXn2B4mNQDRkrH1LtvWuFYR0PpWspU9Q2yLsK7kimerZEsIqEoM
4HwQwzSen+vI10qBtJvP0bWptD2SuTDcVoQxx04H7RYY7rooK1Nt/X9SIMCWKUe4mk8tPmrmASkS
VIZw2pf0pNHeJU7DLUqiZYD1DsYBz1ms/QP4pdCTzJnI8phlUh3DHpTJeoaq2S8tkVn6UI9kHewW
OAXhmRwObkcu/3gLa458WuQhRqQ2VZkV7DMxwfd2OCEbEqX3TY+MXw7cr2PKkmropUeiQMxgF0jm
X8kd7vcLJ905BzNnvnYOLCBcEppWiT+nAGMmeJW5+mUaXl+D3MFTd80SSgKqM8LMLpgPFSDZWB5l
kav+WZju8Zvl/pbjissIeCB+ycy5erJCoxjKhinsl23089v6F39cYOXmOP+3zCMi/tTKlEqT1Jgg
KYsXVeUKY+NkeSsYODJqaCPpWXTnwiOepUg4bVf6p6XVsLphx2xpfBCf3Fst7qCKmY7AE2V2hyp4
GypNaT3bKOda0jqZFMq70LbL4QaNqFCGCQjllARg7jZMTT/3Ac3PJurosMRUGzkZjYi9/P2eSp/c
p+bZoJL5Cy0eUi5ekphorga6EhNsvUhaOdmRkF0AS8CDJsnKwRVkwSlhN4jJcs3Sk6PaLHeKENjh
FZWCXfsZsh1SRXqpyxomVqSwjwlrwekmBvUs01KdFfzdpKm+l/LvvqeAY0AYqORV/sQJm69HiC5D
eNyghJtp50uy1zb5zdQpATZJ1E8Z328a977o/ejNlr3lGY2ZJTH1SxDuOWliZvRnqE/s0dN6MoLy
8Mev8gVmEhKa/9qZxBMtu6IdufqGKIJQZqtaLXEohAaYS/a/mGHGb6iJDPbmIKjsRhTrNby9wlxV
PoVFAG9zynZZefLy8X7U44SLFVgu1ZK9MGwqh2eT2l4YV/KaTGx4JOTNjJBUmA25LZdetDXWvVjb
+PN7iUFshye2JinoNiw4E6e/frVTfRTBZAhRTtan7IOgNFfZX8su8xM4oBcVwLNwb2Rfx2/yoiRi
tCOilb0Ywfm9TuOIemgqhoMqH6amjZ9sGlGo3nE094x5plGtmGzm7UFFr1yy4JvoxCFvPnArv9Nc
hiRQNDbtSr+bg+pfFYM2P7G7ghqFJXMI2CzlrO08nvo+uGvINcWZEXUjW2LApxYh2mdIQSnVwydS
xvBaJxCk84wAb8NcbSa2PjlAWWcYxOmTWfjcjtU6f/IwbeW2HpUmSKwBKifBW9EqDXAEGlDPocb9
Jx1gUvZyr81HYo4iS9n3IBc/+ENAoYmRvXICEiZSbUYCkWFM1NL+QrHfIVXHxjJ74b9XgnJYOfo0
+mXVIfh8MZdzySodXAKKQFRYeRqomrs4XHa+fUXVF9BG2K5h9T9At0mIH9ekt7fftLeKYTbcbmi2
wQr7UNrcF4QtO+gNxAUMQkuI2//Pw77IOkov1rWVNAh+0A2Olg89moD9rpi2PaGmAXXt0RFQudFW
WxZLhtm/PngXwmg5Uqt6knxqWCyBUbhMIIAwrlluGZHJSB9P90sdoWHFgdQqzQr75WGANWURXXTm
hSaEbDcFLua/b90xHznn01IstoI5kW5MVKNdH/iSofwwgUjyn6u5Jfi9iJjskzhdyJAIgYf+vI0n
3a7a7nhlN9XffnqNFRMXrflSr9/YX+xzYcA1MbXlEmvCsulCKHOCeTBtHdoZtazi18cjJePk6U74
3V8TV15C5i1GT/KiRCVDjV3eOtSfDl+VtdVS2mwhZN9eRbrwf8fbhLyi32kI3BmV56zR4lhwXT20
aL/jccoQdA6NgOKI78vJ8y8shIplqWrlpGiWaL7r2KwlSni0P1mWb7sQUVM35RJ1WT3Kmcgd77tX
2iZT+VPfck7vc+qZP3qNbhV4NjwK/fPagDLAik022C+PMNW64iBq+ZMYBe1TRLIS1oymbq40O7e0
vRG77xvVN1A0Qy/7fDR8ysnraC1tk8CL8dSSf4mAQZqjwcdEfIIQPaI6saevI68w+mf1u2Lg6Kat
ieb5XCTH2vPxZT9npO8IwPO4SojjA3+0lV0GrIyJKhXbzBbl0J6SlM2+vL6nCGB377bDOKhOXlJv
0mhO5f0i+Ga75BKRKx/qHdHSeQrIUrY3P3lMhy6rxiRn+yH8076C7zhL/slRmBZKZ7jUqA3I6cL/
wJdO/fjh+zpL2VsxAkNGnNCbqprCgO/wlNqQ8oDdLHUfnDjJ7fXI+9TAD0xX1l7D7LHMbpNgRrsm
xTwR8IyxlMzoWZDoUv68jtNh2i4XBFUQ+A4JNd4OMuJ9PSn1wKmTdhLRqm3uMht38P9iT4I24+py
EeNmBsZoMRF2euRlVDzX0ll9mkLVUuOFJq8lF3LcO4m7VFmqNqQ/uBmnLELMrTSCZVG3A/4oFFo5
iCtEr1A6zn9zpHrqtFC1/zdS5xxthJK4vfOBTKa5UllfZOsaP74rya5xLja+fGpuyT+nLCeGLZRk
I2zenpwC4NB39r5kMfYmFFuEt+3rDvyAmqggYGe1FTU9gV3Dny8l593OgIgnyR++wLlrLNk9s35A
jWhALwHkuYCHvPEb1BiiEPFfpe4HOKgV9f41Hgv/YHxDNx9Yh864wgE+MQw9dkHhN15cmjbvXK7J
tD9tI7pXoarHTcUrumyFQZ2RMcPsQr7C+Ku2I5qh2GCZHF8wdSpK4D2/sHmsRzn4+lSir2JpgTdH
b8Wf3L8utmNAliviht1RQBlJGh/pE24EObfQ/uRxLCEIg5WCxD23U2/RNQINSsSAELewmmo2YifR
XGp7XXGDRQaj17gRzBRlPiavv4ENUrPcXwKOUq6KG3HGSl7/JsqMFp4Y7k/5dIaY82RWvZ971I+F
Iht2/CZ4PF8BIyHxMC9EdXDYwf8d5+vL7eaMPGBu5/J9gfJrdBmf4KZg/4PT/uDGY9iGsYy8c7YW
ejU1swERZdCn14wDY+RfCjgX4EtwP8B+hkzbuEAaZOPwv3nVpHwamv6oItUwXuWCmtICcjs2JXp8
lmCPiLw8+tKh/5QW2em9yWuspiIcLRMA2SlmkZjp5b1wtX8yPTf26272ISfw2LASKP1jejw8FaT5
j1pmOBgyOrxNT9ml126eLovLGZMvDju4uq3XKQ7bEacopnsD7c3hWzhxQAWKM+pFSAGAv4278GtD
i/oeOLeb7e20iTMVXbv7sU0HLERI33IOdsXS6gEh2F5cOmCp6W+m/WO294JNxnFQ7sTfIBdXy5u6
8OmjugzZDV7j5PFHTVxik+lSubvJOs7WHmGBvlo5DCL9mzzt5wZeSBy9BSWj+yT+9BV9YZ0JM1iL
tFWhkVXoZyz70ISFeZMWDVobJKPkCbVPTr8No0XqfwgZNwAsO9fMZaxWL3oO6T/EPg+yja+XSOCa
/GaN6eo/S3Vh9Zn2VPjzBJwvKNc5dH2tbTFCuJCpU/5+RNw8jWW1QAcQ0QE/EK5kR74qYCs9xJ8r
w4/7ZzFxCWffoqPDLzZN16Kwh4TO+mTwOTcSdw18Rj78XBBzJdmZkNkbDVHFtnLCCtUq9igBD7Ap
MSaeZPMBkNxGRrMUNZ2/dWOKgv1iXCZIqcWLZEM/J0k9c7vCZg7ohxhtj7kIb04nnMKuBCFPnegs
wsAw8rHJj8qT6ffWphL7s4KLisMyoQ9cWhX3f+NOkxdhDENuWjIxIxx5rOU/WH4iacV7uW/m+Dam
x2/rd6/Mdur8dIZRQhGV8Sw7V2qWCZo8cERdVKkRaf47GNnHBVuB6zB8ASLcN/wF8IquV+0D0MR2
5o5tyLZj8ZJsCScDqfrUrHSotg9sxHsZF7dLpfM+2yotn1PwfGl88D1jhS3DPfiNwRDLTXmx9FGP
mn57tle+LgdsxJE7IHqqke/YQbEqI+hYykL8LWv7TxioV8tf6/8/muDcwNbi7/s43ztqEtwKTPvf
OPf8fy1RojyWK/w3DD2FyE4EPQqQVhki4XcIhOLz3ummmIvTltdXYXPTFTT6Qgsl9kxwpDvJQGwX
IbsCXf11NqAx1QXOr15SD+hdvyxBLrl+j2rCx2P8tRlob0zdzCDlfsfSDBfBnG8QUdhO4HEHEOz3
nwuCImOy9UeTITVLf8ifWmuRh1dUgcDpXnKWH7C7QCB5uEGWUJLUNrasqjl/fi3QdQGQNqcCjMhk
2AZd38Tx8MEYL1q50rSNdoFpLJkXf65K2+//3uwdlQm8AOstSY7Wyc8FzlAwZP0pM6Sv6IcZBuam
y0kRUSl3mA6CV/HgURKbSoUfD8+M5lL+9eaRogrXXYomgByAy0D7D3D71Avx9OFua60c65DF3JO9
vUT7DI115wcXuR8kzEqH+jND2D8HHvL8fE+fZGGciy5NLOQ3T4MXA5RQV8deWpz1gRtLRXoZKanA
gqgmG47vcMVpjMD8Z9WGbQKIqL0OVb3qVZXDtgz1u0ok3LoiOS31nJdFycx5iAfARFJdb3cGBqSz
pBvbKg4UE1u20lVguuVrrEYx1yZk20T8+ZjZhn4UEFwm0tKdA2tmfRsaJIYYPftgMAsfvrMOUiTw
NG077N4N+oVVR3IzPeOCRS4VhjY4GDlU8cmIrC9DgeLWeNvxrhu+Y6f1uXgiTKyLDJVB858tP0fQ
SOKfgbkl8NiG+mtynqDJnw5C6zTShWort4nmd1Miq2Z4GCwXdhnqIlNSMBxu1WKQ7ZT+HzpvhPIA
kkfkjCCREMscbKmWO1etZu+toisHOjfdIBbIrH1F53E4yU4MrPjVwZvSbph7GV/cCmYVkCRL6CEU
xPVFRAilrUEuLrD2a9ELSDBYhIiRMUj/cUcBVFoaPf4k+6oHvLEvABVEL7Vdn7g+rc0YTMsfWQrb
zl09s5hgpalguKEOhh8klb/OS94BIdBuP2jBwXN9nYySu4UuX60obOg9SLDUZUFt1vGTIF/dUn1h
ouv28wQPB+5q+CxUjkPSyC4Di2g4zWz9XgLoIpdAy61VJDoHXUjnif9+YdCZQkayO92rTQaksJvl
veVrH3iCEiDmTIWgK9sAmxAKpBM4oaNiVgKJbguGmc416EfdQbkQ6jDF7FpCwQQy5k3CBbwBb8OK
zngZPp8IyNtSuAki4Yq0AL4iqzn9TyWr8v3U6pIur8LZiBFVAJow/9kDbCq7a9FeY/4qw5SLkFIZ
RIgwNOrPYWpqp9SkSMRPo1yAj2QcfSRspdHiTJUH3TqCH5tZKcPCWrje2gHHSBnRA6YAPgIZrC93
EW/LUB1KMkvKsZ1zdnB9/wr7kv9g2jsKO0SYZPfsIOkvR3C0JH+TfGUFwfhQY8a/XIBTQd0diZsd
numYkim8IQ1zw97w6yJufdf2jow7tgxctuYBONtw56etCje0i6a8COgpOmZYDdjvYCNBvrOJr31C
FT/C789x53lXAJEKXbLOXF0Mo4Gi+YlSB65BXN5CbxN4Uvsb+1MIHoF57TV3o+eCCSlciwU70YLi
hzVsGgqZTI/cxMFMgPZKGQ2Ti2it3BEGcFCW87rDPWIxC77lkl0JyDmNS+PE6ZNJJdLrPTFaPI/a
bZR6J9osfJLabzhxu/gx8MIT63TJI2FDsL4uNty0mGgiV/AfIeHhclGnB2RQJMZCizvyVeEYUtIV
PddmiYF+x3vtoYlvf2+n3v025lgd/Mt2Gbph9GAcX1fWGsrHsrgdx+mK5VJFq6SdyfQCCXOp4yGo
ggjImC8ftA8KRHavmaiz0VUujF4cGXTZAey05jgeDCnxzMXG76HHpf/Y0sBqE66Ant5WB7eG38VK
niiWyhVVRX9lzxntNnmGDwCD/Jk179ak/ar064LGLKyIXWXpCWdc2IVikGRvWDEuQAXMyeRLErPC
CWbEfp2HF4THZqiBBiCBoaUL50pcXvB663h0yzaP9Hh98+7sffZRAvrBskLfybz8JKfqQrVvUAPP
8OyLwGdWxIEN5P5nlHA7Y5/ri0po8+f51NmHlXnurkojZ7DyDaUtuSj2seKnJrfs8h3CpCKne4+8
77Trsp5fwAHACXRNhW3mEBU1xgopokdD2xgZnVJ0/TTVWcckSxxuZ0o/o6uxeyRg0Ylo6fSmjG3v
8a63ztq5iAypieJVH8MYt8BCXiyE9Ooh/kal70IJCc5ck9DmwZR/81IfJ1FMjo6SMtevSZ70PZxb
F6C/mQegyLTdn3hTz+/yTz7W8mbrUd1jfTQwEZgfgaeRkAmPxG7wzpHh/us3+epNjHNAW4fD2M5k
55ECZ3XjHYaWU6kr2JNMLCj+sMK+h8i4OX5TMuEaC9ib063nj9melhETU17atVAW2T/CX6JAS7Dc
OQoO1DEUn070DvOl/1xIbxsdseo5RyG6Swf/0Tr+kSd9SQkNyfmbfgBNBc3xpBGjBIIA6TZRzw5C
I85jrBBB3/J/MbujskY4N5WKpBroY+LXhMlf0wojIODHHkBxPCAdP97pXzmEMO1mtJo1jw2aoNwk
r9JjxhgLYSQhDCELMNGiqlT3OUGG0JDJjIiUo5shNVjtslYf/stA3jbmQVTEv4GeidxQeTTbvIGG
glBvWElCsZgUUtww3rhT7no51nzelw4HD+9C/l9bkpjyGbQCjssKiaNrpx5b27oz0of3p9JovZCF
cHO8HS1fHJmV64lkE7QsiAi55HrFpF9fAIwrkL8UkSSr/fJJkRt5SwCo0zYmJ1o+YWrhX/P2mR2R
o60Wh3QV2A0spHTyyG79K/WocZVZRGp+kR5rOZc8BGxsC0WghQRw6Y7BUlPN0BN3P84+EGHHU17W
zrGdlnC/Byn3SNsTK+EiksyozFglYhkH/IMVuoc7x0CF5denyljEZqEiEP5ZZ4AuxCdyuEbbpRJC
UApBIZZWyvwQSor4Gx0EGj5h2jWgew5HFLqUfkLhPF+deao3VFqn/zXBWC57VQSDE79WajGUVWdJ
bBUJsdOwSvX793jap3psaHgXPEMx+I6gB/o5dON88hrT4AI2znfO8RqHzbxigfT+g5yhwGGe2UM7
2aBI09e2j7eCQz0fDMw+MFGztMvoVWDzP4bgIGgHafTkauPNEclxS9yS86oC0juVBMaFMKT5Mov3
RrQn7jdCpoCGqHYFyNy+fk6R9ayp38Au/2WKy4cKH8/dJ61sZ0/APGIe+/caJW35ZZ6LbvnNv25B
tCwFtXpI0Et8l2xIRnnk6VCPr3L1caMZSNeWyxNEpBCbQoJNz1OgbGEAKZCOAersTP3o9RnCpgIp
vWGk6rEFe+qmA5HV+AiJy1i5Bq7O33nLMD5VUwKNW2LtHPe0gYHgwM6UnlAlcBhVqt9+gxZGodoK
ah2Bx1ob8ZpyagUOJLuLy5uG8btQf+CqIiVNC50Dmd+8IG1U/UIfS/cUuoL7g0dk09wm0/nZulQS
JL0PUFPTWi35pDltvZmPNIdCIRxuy+oY6pTnknCR17bNJXH0sbFy1up53XNWJPs/cEqWZX9Oh5mU
QMkCnvDExCFJMX6eGwtbJSGQ7gXiEYxgQyTGlJfIRb7fqq4xVZ6W39jjb/Yil+m2X3OaoSxTlbjM
P3Zgry2r3VUWwUPzg3SDnLuP1Z9WTewrBXPtXKeMlrVP4rRR4fBVnH4XeOY/6ldeZT6nVYQefoZy
BcREH8iJpyoh1qQvprjdOGd9s7+OW76B+txswceLpQDBW45CrXtYsICdwyNlmfnIc3eKKSEZFPL5
RagEbM0QzNn1PQ+2KRn+lQcz9sUuHbeanbyobwDlYoYBAM99Z+izjaqv0Vb695trpXGq2nrKZw57
3BT8ix/fQ6yHIeICIoyJWG/mSpSqYW6Uu1GMhfPpZq195WPObQIHguJMhDq2z6zHD5i+9Qg/piRc
SBA8mCpx97K39jnxb9m3BwMsPBKUrCr6ySyjTiPQZzWBOKvk+dI2XGi6LqhouihHBwkOQMjadKLM
J0OoJSZGSeJEIdvqT4YWtkbiLWqOaYmdWFEumOijfYlKJDx+nRTEXyLlr7rN6/Tb3Wa26wMPG7qK
MGJuI2ksUqgwjohbzcazk0DQrlXMYyzTTyQNaB0rzxZISqPup0nFXmRs2lHPXTp8/8YSJBGmD0ln
fbmA6Zs0ExIeeAjkWWIRR6Jp/F1lmc7JNyP9pYVISXHF1lleW8JbjCRxK43i2d93OfvUL1wq+L6Q
41adbrtvMmp6ujPdTHiznnlsIvUmPx3JtKaoK3poxawKZG0FXfOKxfXlUZaRBVIpBLvEiYyqG20s
Lz7XO+xwbuAJRwVh08zNS66Snf8i51P8VIVGEtUEHecSwVCgNUT/ppP96OFrMw/dcDMXscCv3zhd
itfOkIXpK59dG39gk7Mvq+Q+hseHw3JYWhSWdt5FJPCxU8hKrhIcOu4QB1MTCFGkD8O1sXI2D1JR
BMa5qRuhrXWz/tYXZJZTr8MeNwIJ98EkD1+YQV2lPfz0H0mH/X5CnXpNghl7e3NHDBWwEI5NH7mJ
Yg7j5ALMhKiWoWOnApuujdvs0NRwHgLbPieQ3ZZ/JNGcyaw6MtWlm1ftLIUkkBTHB+S58MMFOABt
a/ec79iT9KdnrP7j8ljp3dR7/MD9aBHyhW9CWNAczLj+gSGVkmN5hmmaULPW07axNJ6m/ybiQXAG
M6iPZ0zkzvfPtzkfm8gyeppsrMANycs359uprO7KCIZr+fXDh8EFAF58X/NHM3lkEG4DvM3g7p7B
bobA9TZRh8YgSlfpWSdSOlBHlpYzMWxyFdx7eqMFFy8ZmUYgJDxeP4O29gtRdrkiw55HqNxzS9Lv
ngu3OMQiOSJLa7tCC8+G3aFsy5Ox2fluHfTr6CUmX9QqkQ9fhsVC6zVFJwJA7jUtr0TwY2gjRfJv
zPuLnvD/5QJ3D3JQJquSelp/7/9SEU6lq7LA3hhBJNv3hC5/v5Rq1xl2dFnh430n/HlIQhd0fWRw
dD7K+U+BPKrXbfj1iC8Sa7KD+CPRzd/KxJ7unbB+qW8/fIaV5ewnVapjw3RO7DIWLTMMNxT76eu4
IyzbC0UgUGIjQa/GDWTuyYrBjqgiJLJmOdgCPuropfwJaT2Ao3wKFNJZqirQnfcfG88zl3btfNAO
UwieyVNf/Y2rSFcXehiNlTX3kSmL/55cAmivhDeG6uYQPogG5r87zNQmZ36EX5Ape9pt9oeL6eCa
K2dBasRdpuFQq5jfIcZ85Wh5Km46ri/HOKB/uvfwS5lATt7YjiBaKqWokNCiHpt5Iwd+DzQLnvCB
u3HesfShKpnAXioM1oH319/BOBRZH3APj/TmPmEg7OHiQcbpGh2NNXCHcTua967fAvV4YitzbWtk
FUe6AMjQ87uidpavsdUWAm8R5IfL6SLxkoBRWWbH/Pr3ynkVFZrbFqSF0twtXoyJ7s0Lqz06KJOh
IoA/nkF2kAJThyyOb41+xbRdj+JE5c3Kmer2zoG3l8JXqWzWr4rmzIfPYeyYHHprvE0t4LR69ELl
40+DP8gMlfWXVovEadymMrN4xN2/RnM74C3MnhOHz4Zhcs4MuAoHtG/4Dlnrw8YuSOeRbthWIaXM
S/YJsgieEyGYTVqrSWpBfne3iTmg95/Fe1AVagp9se/7dLzG2YruWYWMk5MeDAR8OjKfHK6f9BR9
vU34wcOU1Yz29i9woG8uaevgZUkUWEmefiZ1iZdUUpLyZIQ6rdh3DYHSwjOROfM3Pi9RX+SvW2s+
HvroKluHnGac7XRPjy8LOwkGzHPeEppXW7IiQQFmHxYA7BTnTYeIWvXsQrhjcMdqdPf0dOa2C4x1
DNsG01R6bzgbEJEvqgpfSAyQD8wsuHSuXj91wKlv1JTwVjeZYZvTZpxI3N5Bwostl61PuAWUNeS7
HRyLTnHmY7aBKthLjoHd5ffoeueb/+gKppkoER3Lr9ZQYKHZrJ5i64TVETaFYly85NQ+CTfyok53
nbgyJ9Ef1D1NrMX0jJVNVIHkRp6LdfqpRebpj7PEr9UAcalpS2efgcmaMnhuSPTn9tdKNqUhp8Mj
UkSlUO6NOmOeY82a07c8M96dFdBMRkpodbcoupNc+sVdanCgNS5LaYdRirCpq6PP88LG0VAfyxG3
Du4JDiBgunu0ZvIOwGraf6XsyLpzjp5UMA1MhJpeKgOzgmOiHBsUmPCGJwgehoXatX+UapnFqc1P
r0JTKsnNdsHbd15gifFBBc3Y+TW5QV2bJsD5zlrxjtNFgRmlSBN+ig18b/L/jbf/Kk3HNajcewx6
pje66Pk2hw9eE93I3Y8tsy/PTkrTYSlR0GshBWlCEXD34qP0aQhWV+L10lv4oOFWwIYfhl1nDxV9
srrJxWmt7vgt7mGPq0Cb/aiFbisDQEPzv4VQfJX3gh79l5qAtSo4XNV+AG8SIVSCzmAf81+Pel8D
dTG24ga4M9gyTcVB/vPP3cUzjvPXq5FzOpV6efsl15VD8MnXlFiThBDj2VzmYoCtCDoXuzi2Bkp1
IJ4bybctGYSvKFhxW3kFsiur0mOVs9agLGvkuoeipT0ubla0XoI4WejBoGu57Kbxs+SSu7+xLK72
V3rBxQPEGrXzmXYGBaUoM8vIvzOKuA9YSMF7Ms+gPaPTWuGHueMk5yOOZ7TCz+ZUbhBF7uXi8ys3
SVlylsHFApANmSpUP+Mz23wphp4BDE05y969fm8JVjvlxW7sf1CjVDarl2tWlpqdbZPsqCXOzvSV
19KsJYUZxEOr8nC8S6U1MDi1x4E8MmhkY+4Qq73s3I7CDSpMPjLy3Z7KbbZtV/vyoGOEBW/ATP+j
M2aakEn0IPmtSXBxyTyLp6/yK97uSZuaXlepesRM4TDUXM4dWX3zd3lgvpWgKQmpevesCjD4lLP9
61xHI6rLJKYdr4Z06AezmSa6YBpviovg5oB9+mHY9C5oqoW/28RwPoEffzxQgmN1dBI3L4orGWuo
0zDkQruFuUqpDGkX1uq2nveCUlMQs9sHEgCT+riLEN827tduWf9XlTmr2eEUM0YbubjMpeosvVnV
eN1QXzrt0b6ts6xYKSRrubpIFpcmdrY6sojU79qFeAfy3+cJpBubEqAYAvAk52TMxpx/3zzZBKUh
lJywXVFSJ3UzoR6XxZixUiRWJBa0u0ieSweeDInDvcYerPdBuzh03l+vv2YP7LeDUT+Japh72rR2
emsBjl6sLB8AbYdqiVeA7amluz0a8OT611EMj4lrwVjaY7CmDqEXjqwrfSehEn6TA2YVsP56ZgLu
8HjW9KfqOvUAwVxGK8W0/dRMS81Y7IE5WmkVufwacq1UMJpdcUzsIlaCBtNHRPxJZS/FJYmNIWUP
hf06DyQ+lczg1ul4l98Ifez6XndLSa3kOjHwqELZ30zxRgXUc0b7fBOIzHQT6vnFdU8oUe/HEyQf
TcVmRabj4MKovHfv5UnbHFgRcSXNu6MV58ZuEFGoJRKfJsk+NMkZ+8BbE1+0+QHCTC/MekLA12/s
rCHLXvdLgxtXQNaIflbtGsikbMkuAekMsJHG05Svmn4LWC+5y6rDna8XISpbyVfWkloCK+ukbmQr
wJeyaXECPblkoVLPNiHXAS4F1CqikDXmabV6POCKrpdKM+1GrdyVpFM78CdoEUPLHoA0iIF45ftq
1WgjrQgqcYJ5mE76R06bl3DKLptK2SSd0e8e6Lg3X1iDd9SDWfSQa6uH26f7qKvDUwQNwcavjipl
baIUVJhEmTC0JwvCOZszmNAvEBZR8Lm8hehNarmLv9EbKCI5Z07NDkBDaSUVJU7Fz/zOhrZ6athY
zGFv04fr/YCd5eUb2Q0OQbisxGh86Or0tOtDI0ZtEKH8tyZS8VHvABy8/1TSNnBqDtzskbMQl4rr
VTjxjvmOYSO20ulfPOur6xVTyS6k7FOmou6KFfSVxw6fO4KG1U0SKPwMdtPJ9/RYIb2j8gow30FE
fshymh4YYx8PRjLrIX3/EXNI4E+VpUtVKZMhzDmLrImeeceJd9pY67Mkrfbtb2DBR/M18WpOOPZN
MHHAoGrhi1sPTNKVPunIs89WYpGNfeFf/TEm4242Kwr3MtFQqvT0YWC1eQu6wPz9we4nAxiDANSt
boxhlJBWdy2EgVz6Rk+c7kZIgVnbiCFXd+kydOAxDD0B/AVC831xCjOsxQcCovAsyUh5/KqRUfUP
lf4F6tZ9+1Ozh9lHnq4iyg3ErM7oOuOSi9hpLqnNUpo2iD8EbR+PMk7PlrqGXBp3zJtqNb4Mkbod
KMruWsfXmGCBAhD1/DuHKT8LibrbgncNQHN4s/9UrlgDaYEIIvZ827/fAFTdDef84qBvDtAKOZ5c
oSLOyjInanjpO76hoOpl5NdSXk2Mfd78nWbIEey0nRphnrGw399/rEiHIVYKBBJVOF9gsfY6GkXF
OE63OnHleXkz0fHJW9fRffp2T8LPILx5k85VhxMa48Xkz504mEQhjHM3a4eL2TbvgHvoWnl6Tyrw
BpINK1M8kh0ecaXke8TW9u/2k08neupCtNL/SIAYJq4NN7EFA/xUdnTmXx4NdpSvds30Pg9Je4FF
LhR8ZDxfKR198ebLf1uLCMDu3VAOgYmZ1Ll1HY/S9y8tHAH/880ADD3KjFoKhbFDi396qzsjTrcl
AJgx2LCfsAAjnpEHVLvKsnZVe8te7pLj4UeSR28FdyhvJ/UP72YFp2jch3lO8gk5xcOXviqZ4/kD
1twvT6sAl/lBJhBZEwcsWdWyKQ6CmxI5i1aIWmR1P424ug7FchN5AxBwT1eHHSKAmRiLoqtFKU25
1hcpOA80klhJE8B43B5OyCvjjPqZl4buYY3AbTQQeQiZnv758Qk0tnZh4iwignOeO5BJ6BUkYCNH
6qBFoBDCDOw+VOEL7UrqQevjbxsb1YnR8gT/oHqN/h5x4D3NyyGrI8T7dyFfpSW06YDpdkVKgZoa
3ThQ9Bd/d9JrkgHwqWHOd7EOtWv/D6DZQX0RF+qW9O+d9mszpHVDg7tmRsT5yfpt7jTPrJUe3KkW
ikAcj25lSet+2q9wUFiiK8xmf4cXnJIBg4YxMPE38rAxJ1R52C3XivEpyvCeu3YAcJQv2MjPjLYY
LyHxFt+RRiKQ3yoLDAPn/8e6pQVjZq0xuy0llPh7X8G94q7MqbGBPuCO46Vxpco8m1RpEJFuvKoo
LFos00cKAPN4YBwchnzBVoWa87NdtPnEZ9P7HY/RrOjojZaPYhqncmnM5LIap+d48DTPobjjzhCZ
cc8vULCxY95TtqB7ZqWsyp4Xeeg3PcuwnVT08yw+kP9/bOSHQGV6bBQCHyi2d/IcrfE1noUSK0vP
6rHC2GkQDFmHm2ShR6CvvsLo9hJAdnGZHA4s7pNM8IJtyZymI7I5eOOl74rUFN3qtbiIJMLki9LA
VClWzzln7x3iwwar9Gtg2L3WGwvMRB/OUAyJylbh+La+Ym961KtVeClI7xYwCQvd7X5pmWI7H2m4
9Kxm9PyyEPhlH7S+jyAmzwlbgKUDX4bycgWa5Zr6u1WXsTxoH2s836wAXCQQCPEXkiRG8Fhg1EgX
bky+556GvTKctYUnnEETgeZFTqi8MlvPT5RBul7zZPOgohpCmkF6Epg+8vayacJaEWn7HSp7rjkM
08/8HCP+kKzhD69vaLcEs8mp4zHBejQVA1EW6P0jgR72YMkyHXj6Up7X/aSKxxaOwJKP/EsIpAKo
0LswxQd30hp0ZuTRSduZXb4KfnjKoORr9vGIHnchzutWUW1wd2RiO3Lo1xyBSeTgqzF3pcHmWGNU
xKeEkEOXFFVeHEwGOOA2Y/Rwux9qclIyD6FTtxvt7SUzw2Yc2G+XBP/toWzFukEHJ4aG0qoXVGIM
bFhW5Ec9RWabUM3w0gNiXl8US1WGQF93tEk/KRuRM2dO16yDc3TG7Rt0Jgx91FqNFDpgD0PVPHOo
e9C7eg05XBtNAF6mpwc4qcKQ4eZ7lt1waJb5KdPJQUGSIJkUlquWNpfU9Vg9B4FWryErLKlK4PNj
bbGmB+O2eDM6At2XEKQgQUVHgQG6bFt8aXTrRTEgOZ6pCU+Cn282V2x+OPX3M4qQATi8EYD27Mt5
QoLBvMIwTqwHpyFMXUr2Er6VKdnWSGxy3VGrdHVDhfZBZ9efK402WJLc+bv8/mdMy7JAOcurxK94
Xr+IaWl0F89GGtwr76rSpC/dhDORXICCDaofbtzp0Jgdxv66AX/QObsSatZK7ELEt7hWz2IeOQc7
IIPQyB60oXjU9wisIuR9R53VCIVuaM0HpwmYNkWq01DgkBpaL/QgzOhVzY8lOKTsHxuZlraeWurZ
a9z4001LR75gwdfB2/rQwbFeMlux7D9Ku2Vn4/eN3Pzh/yUbDtoVXFgclULHPmA25mBHWAFiOb/y
gmnPgkiln+MWTHCk1v8vrj9Mn58c+UDOJbaaDdWOkGmbrbWCXzAuWe0GH6bsC0Ku1SMODnKOfKSW
gHuXfXnO0UIHZUCfVcYiRulpMxXubegsN5XpuDP8qSgPNjf0B5Qdvy69LDz7hFEUhWCt6hrxYpyn
JyLBbIb/XZ1YhmfqLa+iJOcYawIPE6q79GbyziArdm3Tik46e4KzbUq3OpRxP+F02QLhdvNROmq/
QPvASa8wWRj+HnCbDZoaXKxR4fifeJ7iitdj1O3v9NKJvCm58BLTHmjfJ/VG6JjZWggm5M7EhfLE
5c70zm2iAuy3LUaY89UCml8ydT8kiprefEvgylRKXxTba+Blbnhil+g20BWOl2k9gcOSvXvZPeZK
Nokiw1cAgRo+GW4Ya2JHeLbVFaPppdCnGry0IW6Ho+KhakxEEQBCmPz8YPkfNcv4VXA6ti05E92a
ry14/FphgbfCVvtVEOdPnC9A5cVhr9plR3vwCqkGgEg9dHdEP6mypu8JvAqkVz/IuNNbLAqPRV9P
CrFTfsIbafLiKqch7Jx6Lkezmntv4MfOpwqP3rK1tOZLUN3xCqAjBD/V9ETywtVR7WUbGkxUznbm
FbNkD846TH9D3cV9INVh4cqTEbvX9z/MwXLHXqYVWL+5nCiBH+u725wTOWU8e+OO6tU1Y+koP10s
7Fynf8Sc8KuNfaXDTzZo94V0v16KfssbToZjBj+GBAJNlilpTNdggh5ptFfHTUmzU5qF7KDV5YX/
/K30qlBJrF0Rl8HCYY4fkZZDf/yWwxv8MrFmLBjZmDF7DcyzJcgbGiiK2SCxdSFi/p5i82dM8Buu
LgTalz9O9OvBfkl2LB5Ij4mjarjpEHWFfCKAJ7ROgUuWgXzpXIuMiuGaJWgJbwQZJ1qqPloJ2a+v
0u2/w8muPmNVrwQiB8HaBXtnIqnJDv6fqtes12c8vtiI7kGlhcHyg+L8n2d7RM4d+Vg3DaJuIoXc
R+cSNgTrZudalqyhB0ytjvpXpd9HsumNvs5p0XSXwXmJgiip0AJFTvMV2wFoLQPa6e3Zb50nd/XY
Fu20D3sqPdDl2t4C3OUIar2xDf51C9q7WZ2TvMVVaEoR4mxdkUiTiOO8KE/nXd+VTYWL8uuobrO8
nDjte7KFYSVsAMTRk4hK19InYXFZqTPb1ma3PPvqw9l4HGuBdJi72qE8HAxVdPbKheubXUqvhQ65
ncp/GH5YX2Ky2vsmNCXpSRxNdIqy7cwNr9y5Dx7lBMAKejbbfYKu0TJJ6cMV/eIbV40UsZKWdX+v
aRR27rPflTVgsloivd2aFLYjOGvmGjX1NsM/qeYV+r3lLBkRIA4cJ9fI+C4rGpAXpAbaoqxsgyRN
xViXhBV3lL9h1SFqMtOJYBZA6yQfGGW9Z8h2fJBwPGDuExJkk7QA4KHsg0zc1b0djiUtbLnwttrm
kK3ui+UcNCG8uTHUioJdLfeWovKJ20qtHYdHG9ljeqr5p6RC/MsnI28mJh9HoY9oEQ05SegIplif
zWT31S4eCWaxeS6J6mAsUXWhYLojRS8Oih4NCoEKpyKm3jrtfWCLhyu+raxlkQRwjVsPutVy7GVm
QeYiFJwgns4XEY0TrEFKGk4SJiQJ+bnEmyVmQ1bqHsBEY3a0MJ8juDVmXyTeHvxNfuKeAI2dRu8U
vbGq++Zhlkqc9FFrE5cGM2pX8Ps5OwxEXYbcC9dh0WTBxAUl+6dg/sb+qWBHfAc+ZRbVbM00sj7B
hqFM8vtxVThDxQNA4lQkRoVDUVnWbPdKvCzN9qZSJ74MKFCwqe9T4U1XF1gEmXoCjLbyDhgBRdsq
1pUEqXfAgSwX0o/TLptVjZ94pOZHPCHoLXhk/zFgmayARtM4iMZx5KJPgJ2tvAheKkHHgfrnPaj3
hLw0u+tNQCx0SEC3SBvkPYvDU071EwtOl/0QP+8HQ5VResWJPXy9fJw4HlGZAmMCekZEu8Yuavtt
a71pTOqmn07ohQ4OIYMxzA8mtOX+W/nstIsL+DqO5YFleV7Ipr+sysbSyfkdW8cRlzxRkviEf8nc
73EQgCjIW3i9wMWWvB6Edk1oZXps8n7Rz1tof+MBxMqUtQuDLU0ZJdB4mHHN2tpPiZ1BNiKwwC/k
7xOC3WGJp759Z1Btl1kQOvdsvyDptJCbC5meSH0uJSgp5KKWHL4V8xOfkJIMXiwImSmWp+0xG5Dw
nqi5xYKic2ZM1sY0pvToAJ5IfqYmKB/EVdLdFSTsrBp5Fgu8ZDkbgR77DDs9ReKbZhW+F3aqMRH2
qfZlimOqjLCGiiJiJedAuv+1abVUhjZAqlwfWPksWJ3JFiZgEifMPsBi5HSGDMPje+n2pK+OJ3Km
YDM5wfgXGZo6pszfQl1G9A4kiM0B+URRHqFDXrTMEDktHmOmOkcxovGrdtbQgaBvRzZc2nS1Li1K
4PFk/VMgiwv2NXdUp2E4UqPLjtTUVFxTh1A0ZMJNJ2KaE0leqrQDZVdWyen8+yeL80VFZi9BI07h
HyzVZ64wnMBxsgBEMSJK/jEYTXDiI577oLNpVXYThU3I1s9B3PQuqaphqFnnsKsbj5CvVYQ1VX8q
qwoXQWwc4aAhSoiIY741XYQMT+ew8Wjypg4Q18J/S4NWMV5GKI+OCLYjLexFBCl2fyUI9JznXc1z
TJF8VRW73COydZqpM2E8iAyKb/WKXW8724shvVDnvhFtxkcWYBe4W+KEFH3C/DjaOf7eRqR1PydO
bxAQ+45HK2QeoORG1fYBVueSbzRCiqpg2IQVSP5SApxiqs/9EepStaG3BkXJyGzRhKuqOkmx//8D
XTxBaKmpFeotNybleZVMT+/g00h+/ayvhclqGSweqhCIezfIib4yxgkTnSaIHN260HH92eKlqVUf
GTCc1Q9iv6/tfeNvlagVWq42w6RII5/SAYlZg4DQi6pUleF3gQGKiWBdMvSDfD28tGVmTuwiEbA5
L4HVhUFOLgcLMfc1Q4GHAR54WOCRfyKZmffP9YS5i8czUbPAW2Obd5Ppla53jYmYcbk0KaUThpDQ
obpIfEDNcTe/4mI/Xv7tS/2V9i33jGQ6NDw24qiE6Ri4Q3j7AZT8XYKGawMvMwBXs5QZLXHXwr1R
Cz67EiRyZhur5p3IVcAtbUsb3u1UQBDTmVbq2MfFU3Ns/xy1uvisQ7hDwWWmFZlXWgrrL4TXjMoU
2gw2pLjuqHPcJeQT2tPxoOigS+cIjLlJMBzmmUs1oc65ZtZbcKwbkermTQ3l7GAzQY8fcnlv7bH1
4e3CdJnfWAkyzt4L0z4QEbNl0EaZtpj23duaoVfKOW1CQ0Nm1UxdDJNssCZ+8SjK8RDg2ZLOrWGD
xDLOv8KrZduWQSiayEGxpfBLjsvAvuZnv0xwFJ9UI99f6lS7gRjgZfssj4g6f+OYULil9ftlev1v
PVvBNYW4v0dwv5Ykc6UEvpneN6Auhky1GyGlA+hs6MP0Oty/rCCcQpxpnzXjs+/TL619QywXZwxC
2IbyLzoni829Hgk6wzkoNP8da1XfMdNUT6ljWEkhICeiUTkiIuzi8mAHAIiAlCib6cNFN7MI2b2+
U2pqPsX3+0IU40QJsiZl6MN7pcQUKqGCapJm0grlXWyMgyYxyDVklzD88UlCRz7Wc1hZYXnhAJzA
Kp5A4Bi/ypOJTOpsLAP/Enm+hurxvKrFzdxqy48xyPFfyPnX9/ruiTYSiiVRwAqye9k/1iIcFdj6
mm+Y9piQrV7Xj4JsgtjDxUo1H7C5wsV9hscg6WEr9Yz0jMqiX04cR9UNO5lVdHOMRon3wu3hfskG
3cLO//sepZukHaQyGd3D/kzfV2r7DSmCLScvqgOWUjxAMLLvmYwSKZJIFBIPOLp8+MRqjpBr/bUE
3grgRIwz1+9xV7mbyK6b1DjM6T6g4jsbWMygaKgioaZU1d3/qwyutBN5vJnNCKkTaYtnB8Qn9zab
uViUgZj6B/lXpxlG3CmrtYjj8Ysa5VVt7Bo2Xomp0utwR9WszLSLw4XqaY/vXwk0wGmaJ+8cKTci
fGESDEWFIksKbngg3DcerBNpNv1bYV0SBPweR6ZblMmCaQ+tzbvl5TPS4OzoiqCkJIkq9joUrykw
GJs4wYmqnMuNE143HRfunrOkDH4NKUTpCbw9a/y60kbVoy9G+2wcUXdk6VOSnrrgdjILVEXW2ooX
n712qErmxyyf0wME/yPT3qWQK116ceoSxRlTV3cGpvn2HHk7NHWftc6UaxSmojZWN6zaYUKcleqM
wRtb9cEhBsREN4qk5uXZjNNrfSQuGEUSKA+hhTqnrRghsGGoOzmWVPgexkjvphWv5rlUfxQCpX0v
Bz756SVQkCJL1M6IBMpKG34ML3i/SYF3OCY3On+V2OWeuAlXAvmikg+mFFTV9Corcv4bLxZH3xtH
ToNAcCYXRvAAhjcR6ugfzf85wVqT/9nyBbXc45NEbZJoYR8yqR+rVpcH+L77cdr+5XmirE52jy4r
sy6iyB5jmkbQJLdmORghDgZTNYXijg9NlDhujDE7S9Rb7BIuTc/6CIbYyk4sDKBHDgZSfig0/yLg
2pHy+KBhphFn+3pLWaheY1SEkAN4dDzCGLG3FxXHafoc7HGD6XcOuGg0hhaANbm87bNRA7tiyLGa
J3DPq+d7BzhBjz/Exiup5MQNdz93aVQZhsCoHSbQsEKpqhRmPpy61dpiQZ7mOwzQDsJB2bYYuGzu
o8OJc8dSC6/fuiWceAp+RZWKrfuJuirKvkRFlK6Jw6QOn3m0W78+9XPsfsobU8rmULzfME9PpcdT
KeiIEas6lHvie/6HivjWL4fvaHQv1IBsHSHCZ3zSjquhjbOx/z7UXpldAqUFshFxnoArlSCrWVLu
esmTqnpTe4IEPwudV+eIgKRe8c0tJSWtWj5tgdWVI+5M/ZRT1MbMQsvb9F3gFhGSvTeynz59X/25
ag0GPDyi+TFKuda2+sgU7CTDkXOoEmlNi7J/I7JCmDGwnfCvoAQ31kIg+6J/+VXlXUUU7oSeQrkv
TDn4/o8LzOEI7RTGnBJXpGGrZnk20Mo4cs0hOo9aSsdUgILobNs9soi/A8Ve4/isHxFLxGTfj2DP
n5VEvLeTrLqPNvlO2jLZ3iHzqtlP1Z+JPzqluFfH/ScB+V1rEUYpO1eVh9PCpr/n6xUtGgjJ5hoq
C9UTOBjTJxHadJlfOeBkoRQNTeK8dZvV/u6AgaOSHKlREqiNFHKblPa9y8bYNx+1glK4GY+qJiTL
CyKeQN1WRAELkzJR2Vphy4Q6L9O5orYO1QI508qN3Oz3UA+gnpXoBzq6YzlBVNrOTEa77Y4bEPMz
ZQhaJTvytSKdYuiuazKaskbk67bivvqx4BTMmLprg0Cqm5GhEr4z89yEcgCmmDvLxBevDuiizYEk
Bo9bwEg+YkdE0rpv2tczYlMRn7/bF8Mr61c1KIumaOp6JlUr8OnoorGr9cmJ/pt82YTks5BfSmL/
ZLAoo0ngGcy7ZRtLSI2CdqebllB+2ZtWG3g1+iF+lzpcbih44x8xD5sZRHaALJujN8XhoPZwqwZ2
aZkJX0sjCXDnLY1EpEQkqOTQwmrRgtunyT6JrxoTkhOejRARTMieZGz2f6JYsG3hmw8Rz06fsGjY
Nua4BrUuqCIJTnWj2nsQe5VwgzsVH6WolX9wg5EKWIgXo1yNqRoSMkvMzzcSTOjwMeCAOKIrvAsz
+ES9o4qtRSSpEuvMvomV3t1EQX1IgnTCnTI3Nx8o9+k+RyZzzcg26IUT9jkJHilSBsZ6qOyWmhql
oxTfOJe2Yvlhgduq8Zn5U4fCmx2hik1HyFU1H3BkF/FxC9XcKmWkBop94J3s/jM7aY2AHXxo4/JE
GHc/fk1Hi8eOxlxsZJcYKDMDBKA7irvqiFgySLqEBK+zqTp+x5ckJQVDewLWmC+yy6JecMd/lazy
HIm3RlQt0YQHZDYm8Df6rVRN6vyiGDQChCQSUQTOJ7Ks/SOD47nsoUl+xJH/gSSRu2tSW67OenGM
4k07pTuUAZ7SAVpCvPajJOV3rMqBMGhLMv6as+1Nt4eHJug8sqLDwJYvYnD+9/FKpCHuibtZQ/Ml
GO7OqQuUxzKGb8qhHgPQUCPdt36FhWU80OJR/kvtm1G5j41PQmpYpZxIsaV4xJ3u/vxm/aIgR3Ve
5sroVkXLvE2bisbyvm+hedCY2Q2A2Ahmh4PiOJFbGVfqkjvZbZJJ45m27a+zT5PB4kRlSB/d1E0b
huZTLLcKC2hF0H9VILeHS97ZCinZdVsIv1fI731nOeBhu/woaBdHk5BBs7BjJvMkp1AOPtpaAXwT
mHHgbxkT+g0b/etphYcr1qxL2I+kyrnuHYTu24XOgvWbNE3ZAvApNR7ddmXthl0DCrwOfNi7Lgyy
7SFmOqjnypItexIksK2XPF79U3QsZXedCLUS57cFSGlrj7KZTzMhFGKqB2quuNsVhuqt9Driwn7t
KINoQ7R6BEqdXN/CUIYMhXu/n3aVOKbZ0fGmK+A3otKNxCSeStiheSTJKXSxPFQ4EvlpeB38ONSY
AuWjKITlhZJB3lOYIxvwynVsVf5nkCr1eyf3nu0x+h9HUzpI0kRrdgy3RjaGp2rVf9/7KpbE0MHY
SxwiyoluwO5vM1Cmk9NoB/p+pPybLF2QjX2+zq8rZMwDE02c9J3dDReSUW3AUTGeBdQtcNE/SuqL
E1GUnMf5M7xBsehYXZ9qm9ubEh/ReY9DCaQw/PrNgsjL8OHXDvrl6N8UwPZc4iuA7zm0FapYBrs6
raY/Wuq6LpqaUEzDigRqfoDorHDDnUxaoGhE4PD1BxwCjbnKvGp1VJvA76mDfWuzoW1eReLb5lF+
p/qtCYMTCsgAxlymhacLxr658V4sQQYSh4RjVqg4JNBf+zIkLAxyXLtAtQ7saYi8gB0Thz79+n6z
izwDSy9846hmg57Ra+2UZzdsN5QPoublmuCdWqm84oOPnc99hYuaPBE8aEO5uscw5onl2QuSAO8F
TFMr3ccsVD52EFfFu4u0x/APDtLVxWR+grKdqf0EV+hfsIunaYRXagwR7nhNWpo1b3Gn8cw5yqBx
wvuKZagq7u259ZWIykw1/6Gb88jFO/cWVygvSKiJ0XjuDu5jMYF37wgoEmXJbTFWhyKlSiAE6ALX
H38yKC6D57XBKmKUOXy6kOYa8EV2zRxmZG2Gb21zQq9IzQvEQhKr6PxD08NEUtPQXLcsBgD8Xd8K
pXlvQLuEmCdMuDTe6whe+uaprbY6ckMK36VF3Gyl7whM2bOwWWxmErm2QZQc9ZWwa087gr/FXTE6
fPaScyrDgfpoQBJWaLPTRqtdJn/OjLtkJgJt8DJe5QQx4sW7hnikNk6pi/L4pApIO+WgaRHPAkgd
D/HzbjpmbxSBMY+Vcb+bmoZrgFIgOuz83jaQW7gHjr1MzicpfdVPBCkHGz+funF94o/uvxtlp7+w
Icq8MSpmEb9KdPtRkjWoKhnh1n72iZE3yE6s3pnwYOoANdiQf8dit7Qnv4cYvPDBV3X23r5bZm0t
p5HUSRid8y7Gemh+0iNBLqyC7fe9cqLd6VjAlt6GNTtKdWbPhM2OMYs5YTwGRS2DDNqOVm54t+UF
k8uxGq4cTCKiY33ngzlQ9QNKspgRI9SKi+rdZZov9fuuk6m9I2T2kxn47w8nYJlvWOO1VYylsd9f
bHS5rcTUS8CKvtUHyJMZ2EcuwoGTqdb/4OPoaR7oFIE8Omu0RoNGMK8QM+1T9FFiOAFJpvDx3GC1
w6UEwQttE8WMIo8pCKtHr4s4QcFKzdiLqMPCGqRav6TCkVFVPoPuG/TQHeT30RVZALdtDrNvnkmi
QISsbKpuguzaaQq4w0CIAEWf38bwNSAccUMmNLZHOmv6tRNRctZDHk68G1D1PNfS+YRXnaigs5kk
OcS/HSFvEgJmno/RxYgWYMjcemA/bkS/wLho4s96wUWCQxEQc82oHPAhxxyzpmPM8c3FsPF0u22L
1WOL8YSub4hcemZfmeEppONB9av6oROOGjQuYS1ojecuQCY/+OLBknRU7ZlG8PUag1zmCTGA3oLW
gXlF52HcyAO5GFerCo5DR/25YAmBVkcH7FofJG+G4GMxDUJYqjzi709MIo2W7OgHCkAtMrf2Oihj
y+iW3tU5NdqZEVaVTn0Omjre3qLwhO40YzOnnOLxVB4vG153reM9pH28gkaHO7F7ozCZkxAZCpj7
aaxkqqaPou1zX7lWkYNRArmt88bVoNjv5doRtu08u6Dpd5mlkJb39B1n584BCbRcxKW0VHxKF11G
p5rs8qHtrfBGCMD5vCBJGMP8WSJ/bjlF5HAGde1ma8DUm6XcULeLcw/Rm4RMu4V6sWrlGLIZw2tC
GqtGawPqBVyfKGmqlnyiBep/Flvb/5CtCcMeoyAxYx16Nxg1ZdPYjS2YFInrY7jtBaCPC/osBHyD
FnruWYTR+afcUDogwy8IUiplgxdf2jNyN9Pg+80yLRJDgi/0v8yaJ+MXKXoJSvBmICGUaYvSh8fz
ubXPo8uGZ8PwU1X1AtW8AEfmf0ssegVyPisFLrUnHLeAE2VTeQvS1QJ5ULGvCHzD8nLdNryoRQfU
TJiJpKbe4F/C0eokJsfSrHg3rfXBcmVeUad3wgGqX5d0lBg9sNJytcCFDcrZNIccBpZK4JJAmi4G
3mmmt01pqreFLrRjyzd5HZdJGdXFdIBIwTiwrpIcCujY909FAOEOAtdjHChKHkRgdlANohhFeDHk
iGp0bMjUcJj6ncVhYTO5f3FFC15j8Gg4jAUUtuk/APnWJKw2FS34Q2gAO4tLrvg3UfRPN0CXqOSn
UiIKWpmf5Mjft9ZX8svuSgA5+eM+foLop7seP2mpSFptwRWTAm+9kCUaSclrqmv3BOkE75Apq4+t
ioxOF0GYEJIA0IqEnFvIUYsRdCilJS8tzYbdq94udgFFwnaQSusZQ6WW1t2kncyNPNOYFibxHFnX
dsflBQZmTN6Uf50/js2NzLidD28P9+0ZJYvpEvePWhAdUIO6IgyMDt5esqHT2KZmE7fLMucWFJ3/
ig4piqjns4+Ctex51DK3D0hcnc3p3VKtGGHOpKkV8ImdBbk7TLbzJmfKAK4BnXK4Yj6UcaSN422n
gr1nkHZMnf/mja/UBjkNGPJFJ1LM8Zp0H/rcQtBgQ/ug6qtNI70MXASurYhMNpXyusjPDpCS/b3d
FwZt7Y3g7wjyd22Uh9rb8YRLq6EXvTOKmMKYKVJnQWZEuCpvur8wkJN79Unh/e2Rn6PMhtCaYAj+
E3t8d1eoHXZZvSjMm0BcJHNVUK9BeSHFDucGxKxgchNlRazWRtXIw0mXpVFyKTQ0eRxkWHIdOdIr
n0kb0aLXTxn66Yc5z+qOr/0i51qibXl0po+BIaEpjOie/y7mQE2gvDOoyLI66RFGfad898yZWbEK
Rp7HrWrXRIEbEUzFTMQLbFTHu4iVlP8bF4XmBA84GGInogJ2iiE7JrHijcU44+EPu7Mw3Avmzrh9
IzxtpzZWVrQ9IoDLkylgIpnj0ya2vB7u3PKQE+DlnmtZt0HB7KWUOP4SkjKIAhIN3MCkl3kh07iI
+G3coXFbN6DdhgBuuC8Bacb+lmVVGLwr2lnbLXf3pdxz/bmhY5tvGLOW4Ta3HXJnfxHns4gRpVdQ
Vognuh5gAKW2fJoDqnJFsYF0Gf4lba+QATu6+VvcEgfBnmHEvHdpxTc5QMiRmFlfWt5aJJYvJEx/
Nnt/N58Qj2ldmTPwbJg4GnsxWzL5Oew92sP6kxN5zKvC7dbNqhP5beTnlualFYykEJf5lyKazgKW
efvGmnnv7U7NLThEctlilTtj9sHGs38+EJayOH73mHYYQ+gMHpH3kk34I8hZ4KbqrZI1RnkutH2I
z42y+JtFD3anNdMwQyCVcWDABQ6YpCpHa7C5bpIP12bAbpBCK8VxwU3OtzBiR4LvOdK3k1uWkM8f
5W4GFSTvCjQavnxdF0asaBpohwz+WibaSboe4qH8pTbu8XvbTZhXJTQuHZ/C7chgl8m8fYOqBk+o
7cUbhyBwSTncmEJZdgfsk2Uz9oLA41/yM15vxABcdFxp6JGcI1u/DNVKFMivZLLe3u7IM0RcAb1w
LiST/K2k1oayxenvDAFVaomGVoZzEdxpUjP/Vx9omlYm5YVCgVYAmEFbb65DaJnpHLrcg0e4rS+o
nq01/NhpgtOpR+gL8KD0ICZKaU3s0oGws0lY7pO8nwvOUdU60tjXVX17n5nibJ2IwIYlA+qv+2V/
6bavgaEqAT1VRueDD/Wu6H8k5PCsCnlY8fV2L0S21zMGvMYFJ/3HuZWW7xtg2eBX3Ox1I7+cVH3M
aWgpjm/ABNDEItnPTUbRgdp1JwR/6j4vqdnLB+hvJljcCNJw7hXwiuoOV+VHbhn5Raw8r3sY71KN
QURFEPVPR4OOzE0r9ej2LhzVSG2K54toFxwqcpT4J+wR5/MRtnRutALYdcV4YXw+daTd/cK1u/FL
6liGS0gdqfHPQiY7JjbVD3LT0+MLahZQqB+y9IqoXkNuMviGZpE8MuaUFeczJEebGbtvwugZF2MM
Ht4GozDtj2S1bSWTU4S//p+Zg/oUmDl0EWY+Bemg7AxC77A54/R1RzAi6uRitb7jAWk32/lj6IMv
LjA5yQHFN2gi2ni/XR5kQrw4VfBySzZvAjqPN/qNPw27WSkcPnk023SBtbJKK8Q9rhoIiMHf6cQ/
n+sO0RiWG5+Mrkv62tskI0mcV088PisD7d/urRHP3yk31lZdOnz52yjlEnzwEQobgkBm2A8Z1bCA
/ozVhplGKYWg82CBuSqWWLa2jgIzFEwdm5nf110PAAMLw0Hvl0m3JhMW2oY4yRqyLSThzZlwQTcw
eBwsw1kROztHpdbHjoofTRg67yn42RiqxpwYDIPGoDEsdNB7VnPsyE8886PvAacSDlfRr6KbI2eX
TnjzPqldfeH6ld1pNKuDxqhdQ6byuWRoCrOAn/VKxqjIyr7umS/pDLvJT0+9fqUGazv8Ne7EbODX
z1AD47hMHCRoWTZenyq+OHIJyDiQLl6C3ol0Jrvsi2gnABfcAnPtqJRi7OgDJh9ycz68YZaacvwJ
vef10b7Az8pUrqyfBuTrCRwP5dKRV0razzk71F81cTIqQqbwMNv39OD7Fj5k7Y0/arKc7C701SVD
Id/djBF6zx1ueykGvRLDyAtmJPE3gLAy+mrQFIlhP6NPNhRSsDIamzqOzDTxRVBFQdHaF5HgQAE7
0BrBLjsJaKZFPMMbDKToQW/8ojgjuHLLC6jqPrrZYPFnGevL6MqVOBxDhNHF1kqb2ym00V1FB23q
FvlluUj9u5qW9jCH0jnK8CN1HJD/wcY/bu4//PA4Fgw+sshk2hXg/QPAynh+WcH40QZn3Qkx8bN5
V/JmQmIbeUgDwdHriTvJxSQQXLJzOpNRMLBPLJa1bPM14aoBdCtMAUb90mTWcsx077EXt99wWoXA
o9fBbbtF5rE8QQe2BVEK4UPPwWQkajBoe5vNWMFwCfNifi6w8KGNJdDQgucGnywsneQbfTIh1ocS
EgRVfeXln7vXjc9o2Feza03qLSDdiuppSEr/VcCJ1NXzpaWlYug29iDjRt5CDqx3couGhcOpbPkl
wTe8FzTbZoG6jPomr7I841DjSS/BiFDDGz3LXNERvQBt5uY3sejx8HRM4ac7DGmm+NJF/OubX9V2
ybSMgWpqbuzGi0YskgjsUT2df7oC5xfI9rbYVCa8IzUXMLukHW9iYB4Ia+4yp/CbEiBXAsKDKG/b
VmJI70KU7MR47XSy06oaewsij0S4vBTNo4VLZ8GtfUN1TLhiRheb6ZP/yH2LcF8SQX8GIHiwB9L+
RzDiFqCp3mu55naO0TRhY8ZeeV8MYxw2skZFjBd+6BIYFwR1Kskpl2Yx4QOac9hN9wLFaoRl1IOX
F4121kS5mJNw32X90jHxgqq0pdBbrCfgIttvnzo7oJBmjKK8cscJOfPCcEMVVt4l2cN5NeE2Oc+3
5u6ntBLh+ZnuO4kb6EwoZUvMCipjr2UErrqzavzwjQgke0ne9TFfSRjif0cVlnx7UIwqYPiZs2k/
BtPjfJFUEM4kksIEH+b8JPjsjfeSdEb0RIueGPswxJ3qfIdhqXV3cIg/0NmEIYTqbRk7UVbH3Wz9
rj0BYN+qv1ZYb9j/5RToIiFWZ05XW55rs1BojbApsl43RtKc9e/0tbMA5HKF8GegbWRwxmfhUmaj
w3KfpVx4jAO7RWSC5ELZDWZtDGiXtpIcskBJBGgEBcTMq1aXfbU85jp3WezcWQXSoNW+fC8MequP
ZKUe6LEGKN0bX1gw6qbVZ1PJ029f3+Aql6cQW9CjXZEcdePFQeQ1myRocFs63+76QtTBZ5YiGRfU
8yTE/mt3U3oo6eRa9WyZ+j/Ob7vmXiKa3AhNqZv951mv11zsVSSpdS8U87Q+nBS68hWt7mjyt9hA
GF567AcdwycGNSu2FGts/NxJlXy4j0bynvOqL9bsYDkZojgcyX3ecMROe/6nfbB+PH0x6DJ9W6cQ
u1hX4Jd9uxP9af+uaaZMVqGKSXMWEFw4aVgqfLyFrUpZ+/48odcv+v51+npNXtRu2TZ7seAjBWlm
JCfjQK6BmosmDr36dzVBNGQ9JXCmOqgVKAZO0f/2gyxI/V7aYu2cHf419aUlFhEWCNYaTS7O27sM
WaHcCkVnT+A6FkMXQxfE7P5hkdSYTF+LM+d7xveG4I6+gWMhNvSXiLja5exKqHSisBTzgnhmyOKD
lP066iaA93MvjI7NRiwJvSZ5uSII3s+YAF5HG8K5rq6Eyt5rTLR9EHn4OpXDx1AgUHRgul3h/ZPf
ofcuPsmj6Hqx3RoyFvVcg+6vuubd1eO0MkTWszvYJLQHgy1YPWvhJsfj1O42plzG5G8Pw9+uCObe
YksWzcm7gpyKUBk5F81HgqrOv6gJ0+4KUcpj62R4Ooq9ZXJu/7KX4m23bTCJBOI50YYyya66dJ7h
ekodyH6G9zgqse/DrZE1ANXNJ+BPGdX7uBGJCyMJAsssyZw9QkZTnCCb0eWNdauyvTklJWPUrtak
Ryya5ZO/Irgz62+1viXJVT/yvUr74fkaoSHnpDpeIvKGfVW7/pa1DSfT9hTbhtC+Bb7Ony23beHP
K/o8UxYIei6GB3lm07YzAbJaXvLQUKCIKrv6tlnGCdBAmFQ+c6DFZ4mRUV02IfB2DpH+MFG3K5Y2
1LtoI4dJcGI8DbT7DNbUDv3IMy3cxSX3FotZj9AOC/4ri9cCORomOAs6qs+2upKsLmgH8gXZr423
UILuNnm71v/bMIK8Tilbk3VGR8Djr9YAW/Y/aVcCpFQ6PaIRJDkiz5GYoGv27c8UrCeHfPkF8TVN
ATnc+qFx1cmRGTVvdzEyvzgwjZwcOqcIZjJJ7vvxHcLaStv30sNtF+2QPPmVX7h5tPDcKOvOSJFo
N5Po5dzmLh1UloUM8jcujHcqGQJBC3WVEbZxDR0OIkkXn/1NF8SRc2FiKh8xV495wK/gVZZnARcX
WKGbhP6uIldF62jmFebQOtzeCYoLxZcnTsIFF3EJh1Oj88Mli0snNhypY86SBaGkKjBHrAgn+YfR
dZQ09l4CGqyWLJmegemLxaNZd0CSV4r4OcigAWbnXj3eX/dac1CVhfYM6y+jGbiDHA52hpVURJgn
gHIsnN3JpSGDovWeSqROV8f5fkICcyqpo2yinLg3uJLqEiYt2wzKIaAU5ykyp+23QnBv+Nq/84Wn
1NhDz97M0BgX8RfiGLfyTXuxeEtzhzud103bB+RcnwegyL7u4ynbg08hG5MdbVlESZed54edVh3F
3ZopVTzU6gY2+/Hior8I+OI8/HTcfFPk+NpLDwR3L5JJKJbLTCK9+017aREC7fMI7kEGpCjj9WCG
UdKl6OnTPcE/u/h+V6ZAa0iZjRf4h+VvmTKyc0Rvt2jmSwRUYfHodfs5unuXghUnk2Rw1xOaHd4g
i8bpytz2SeqXgDS0Q6bzssm/RTv4cmrdfxbIjMfkp5B0YC2X8HcSwNo9wrQbM9NWi/4L5pJd72tL
gBCLouud1iDrroH34CT7Y6ykdHMSfAxlMO/qLwFOJKGL8ijhh9VPZPn1zV8IN3NHMW6tZ4m72ATc
Sb4IolagzZ1O+ldlpv54LMxdkbvH71trGJOhIj7yLnxCwMGdCzKN2eJW4BBzeLOO/iQKMl+TItMI
PdVymySfkHtnLqfDWHGZZ8+OUigrt+0WHkezPiKf6me6aOK0ItZddNc7WWTRa2b8Px6xu4w8JiXm
rHqk+k/dy/1VN3e+2n9GcD3y+hvlCDtUblMFCyNbEWr565z0jfZ+BF8gXDGC1DzWrPawn5w1GNRE
0KSyFgxxZlG5TY4qgSV654JSHNZ6EP8Tg+OX/7FjRiGNnBTYcgHnhmZwgMRg36h6ZFpGwmfFyMAh
N5C9pzKsG3f7+xVT2FISV2RqcDItOmjz27QTaAlRIlhPWe23JDnV3Y9lYHqLZ87SB/I1gE4DGoTi
D8WIaE+Hnez9ATgzTfuo6yLnjGEov7YnHZZ1Nc3syKSgqDWD1w2/6DFvFIM5hE2M6xvshhTajOZc
vZTmBlZExO3YpiC7Wp9AIRPX3U3wQhusxNfB2sNZJZjcRbyXEZJ8vd5abhbQqp2h600mau+Xj56F
iIZ3mOqEEBItltMvBbGFfGZ/aGAKqRY8k6tFNKT2nUGtNwwcTWoRUU6UqOktsOqwyhRmk+i+Llcm
PySZyODYM69fZBWUMoUA/fdQA/yF2ex20oS0GbPNhvXomuHoEA1iDjqy9BvMx0wLEMypMFrpGFhv
pt/5KEP8/3JLwhcbmLTD623DyEmSudfS0tgPzUXd3hQFBZwDtsXq8hwPDGs0LScJTu9N7IKeav4d
csGFyDs6RZj7r6cMUc0bnuWW3KONr6ZvsOWCHbUB+qCrTM0uPOeerP6tUod67O+zTf2NVrHUXji3
GBnuOmI9ovIfqRt1iuQ6ufkwPWhyzMb57q1zmldiTf7XHsscBhNOoDvOUY38mcuhskEtFUTlQXxm
hs4wJZQNmHi/VjqtS2vpPT72tImuJcancf32g4P6S7oVGEZBZVZYoJscCmMwTzoyEK6+OoKJCE2c
ZisehYy8xwP8plozfDILbeikugu6pjni0VLZsnQgjHkBZjUoBJzOXYaW5qSjYNm1Kb7p1nziMIYf
rBmITh+SL0YAPsS5z1nlP8KxsoW9mVIWd9OUpsF91/XZYUQ9/j8dAnCht7rG8lP7Fr45BYd/6Pwq
NBOcFgR93IQGVyZDK/WhnQnFZ2tumF613DBiNkfviqiuKyD0y1TF16BW3RE8sEHITtaCOQ9hWgpw
knAt61BdP8pAMt8XPbtQBFHAPmkH9Mez48Au2Fl708G478UaJzsiOTtyXawuvmnsrDyTjCp8+b9/
RU/RifMue4LWkslWpB7vZMcCSpHqp8bDsiIe9QDcjvviRXJV1cOwaOxyPtkxk0ktncsVMSvbxJaX
2MDg7UGQo0uNtFxdkcyYZTjRLBFBkdIV9qUtpqI8ZO/pSTJYk1HHKSSHxiHfIWtGaEJhsju551CB
mTr3Ffsm6PpE6WEvXdnIgrRDg3CnFWH9vU7Y2AjCsfcvZbHBaGD2R/cozg1LfLJzh4Ad7XMVTUvL
eanzNirzTrfaXp8HTwRt0FVbdrktR9xKL//gvv4iVWp1jcGbn+f0OvlJGQydUXSH3Pp+G5+eNd2e
lroCPpAHlznX25GmivLpm2psyQ6k/Ky4KRAgqw3hpPLbuSU5L+c3ww9JniCbn4bkghLcZhwHnru7
zmNNUS5RBP7LE1gdhqJObC1dg1aJg6TC2kOzWhcDfGZPYWdIR7UF0J7KDmv90PfoxKBIf2DcVCUX
Og4yzn3y8urU50Tx6zyxJ3Sd5IhMWDZh/TtODpHncPdRfdrZ/4E9jH5lMi7VN9pSS5Si9ovmAKoS
NdODqkFMCUCHa725feVA56BdSPM4HfHomuwoYTVJHk0vFDzj0sYMxZUfVQT97LmZ6sKbbA2Xz3Vo
6mSp+IY+N3ZupC/FWgnk9j9OMbeH51RedRCJWuFRGJbKj84L5epB6sw1MS6cmaWyl6FVegcXdHHQ
fL+aw+W5t5DW8vWM5XYHfeVJHhZtUJcHSQC+U9/iIpv8OTezwTv/+sh1FAx7zl6g1zTk7vGoWv22
JA/gwxC0zN4LkpbgE7B1ySf0fA/xszHR0MhnjnL7mZi9PLxMMMv3ACTugqQbUqVzKiWTINelVP/s
P8EDCMwtRkacDTsJzTe7P8A+2o36V8rtZpXu6LVoZKGFAUcPqfS2oJpSi76T6utt+/Qx+AlFD4Tw
m4modNbNwApaWHDj8BKsziGH4cIX89yCF3NN7hBneLOvAt8tYWIoAl5iVoTLdP278h1pVa1qnVs/
JzgD4JnAvIpewbDb99YF6g14yg6QsmyNp1Yak9MWTYYjI59XWPFmcFVbD31jxm7s5qts/2pKNQrC
Ey4xMQUQ7tv2fhNo3xe0/njbv1UTjK4YOsMrzDc1L1CTsVdFQ7hpiNZ0AVGTOnhs+iFHstBiQI9Q
+uYQQr2Zn28ypl+Su7iGDCAQ6Pz40osvkZGUu6He60YBeo0jpqAvGB4vOXv7KRdNONaWcHSl6w18
Fa+s8OjDzwr52RDhLLi5WdzXFNkE2KeZfN3lN3vbT4N9WI7GFNhZiNv4HZvUNIFyvlWflLvgemuc
dRCNb4i9ur75aQ9EqeeLejOmzQdv7JfJXOuJd3igzqXeoFqYZpNaVoJcmzYwbSpSnY6938EWz2xy
0eFlm1ArW570eEmy4yz2OM5J35DtVshpzrgT+KO0QnHuvBX8fIB4FXeQEgKnB5b5gbx1F6VhKlxs
GlOd6ozgrVKyfo7B4KUwh9o9ZzWpBgVFK6cNIc4GvkMRY3XmzAdLZiDTPyn//obPjiNjZTfB+cvY
aTDzUlyuIEBwk1lq2XC5vz1OG5lbK/q8I0SZfqdRuutOLHL9MPFG8nV58NkdSMVOMZkfwAWugbYl
MrMDYeYKj3tfuSPBzXVU1Gx5tKtPjQtT3+gbgTbNIzkDZ6i2459nITnE5BtKnwRV6MbwFZ2D1vhA
yNVsJdWiT9J1Hrne2w3FYKt8l0F2eoa1zHFw+XR7JHJhrrnhmPLPgxv/0MCb/5O4W1YxKDkDJ8s1
YO5IIk8hVBcQ+LZd/+HsR2RxdzuLyM9NGugQfflWOtoF8/ALf5xnYs4pmi7DIs46DQgB1uy+mZFZ
zf4gw/iXpyDgH5b1imsfuh1Rxr4ZtV4M7dtqkb19Oqc+e/UubWLLG+k9VR9XaIoTK100wR8u/GQB
U/sP+H3nfJO6q/cRSSV89/Gzm1On8OMoRfxGyJxRfzm4ghkBslQi/57LjjB+C31PYux8rtqmVuvi
TVascfjtvcn3ObkUXP06mf6E51RrhSk0InKaniKIKeH1CPqM6egZz69qQ3PP/eGKh6q5bjeFlV5Q
31wqXrARCLaQzTO6M0YTQITAMLmD2SC1SA7F/zmjGKAMydja3EATejK1mCBNbGyYXi6H0YlMMxX/
BUMVnem3UugK3ggkMZtuDchEIwavykF5ClKYc4DEf4E8rBftCXl/6W/IHwX/QcAWnfHAtlWm4v+v
krJSmKQXCe8Gib7HWPmWqAH93eNsRH5WeD0omhhBTrhoZuLmpDyPswFccmv6q74MUSDF1LDXVrNz
+uEAsEi+ww3Wtd47adWfVCboj56Ii07kPjZm0PPCKXWU5mL7XvfggjQJmcpUDi03pl+1tAR4A/H/
4bXG0PVejb749tWAJYWW79Z8Gr+K9f8ywLTmeFArCl0co3n6RWZKA/MozszHtK7Fp/BPTDiO2/d/
r3f5pueKFk8Jt7aCeq2KsNdRiReMxiFR/TWqyEOo3AT7S9KCqTJTlLKgGOCzDX+PE1IdVju/LzQG
ZRwTteGZVbCfzRMXpwNwZMsdLhWRO3YAPFaRxGOUvaToUQZF//G4I/XaeazZatsm7AwhXQjZBeFP
nnt0rwm2Ab/XD3sOh3XzfcoZ5B0e6U83cLYou4Ze8uigV6QEPI0VZHi9V5mi+Ez0DkRvthrZhrr1
TzUz/pkk1NJkpKHLAIaPZsO2TY2dc3r4aEtESID1cRLfFkWD7ttNMyAuNi8A84Rr53xTaVZAcTyT
Jg6rbSTQyOFUcwzm/GchqsqpNNOqx5RbWgTpflXkp0RVyQRzm3UqskXTAlZourcrTaQ3LgYu2Ccv
MY/HdIOkvyeSAIX1jVdAWmSKJoZZpSaDk1vssMIyZ8MymzuMqXFDMBFMfo/n2W2jofwQzBewyNJQ
ttXdR9Qtqf06zVt2xcc2GabEWnF5Tl3wj4259v37POnEKCPkrD6rw6vwiti1kStyrCnQi1+F4oRv
+1a1cf2Qc3eqrEqbZUObj4y7KNhl8xOs0WoEdVIsh8FsdF7W+jTeKwkHE52mo1Y3xr2ji36ky7iy
6IOLn60X5hqLfJJyEfiGHYS8RP26GqVxkVAlPXpY7CDKNZ0jziqj13iU6++q8HhcZIOH+T3alY7U
LQuLIIDPeSpFS9YhX2DtqL4/3wVlEe1CxrSAscw3TPqvbTOA7EVStEndHLv2bROznHFQV6RK6F7y
h+rkIGB7FHbvybQGK+hHZb7Op9pGGiFgFPmpIXxWiO2ePPFqmDYHPEYh3XxQcAJTij2VdK5TJ4F4
7mcZ73fA7O6n+EQF6JOZJRRwn/kikoKW8+zX9NbOfvxo80HjpXNtpApols0cdxN8+VyydXuayTJ6
6beMOLDICqkz/l6YdzJHfIrccvJXI+habVukjxH7lw1Rn28oPX9lN0Is6BAq5f6jZ9lg+4vfiy9c
Y66lsbsgf1qvJl6m3+83Z/NXUjsEtSwj3dwfh5tR7p+Vz9OzNn+XcXuZM9RShJ0o9CsbFMU+JgDR
oPoOe/KCruc3qrkQVcjtN3ZiyPz93lEiDciz7fVkTwCibJx+5lIbB9IVbRG7+z7pT3d//qTBtfxn
orl/uCOjXGhgHj8VkDOEssnCaF7LeyVf/Ow4RJamY5YYBEhlhDl7dObqNwjgdZeT8LYT2FN/fPpd
d3p9rk9OraGNTiKdv2m8WHFYol0BCoPb1fBcK8D+u3df2krhNebZpGSiXjLEszetFp15Sv/6RAXb
KIy57XLL8dBzHxYstttpgx1CT/GdNVNPbPGOPBLKLM/e0gwo5Xc53ic5FPsnX//DsIZ4IN4b0Oq7
USSrwtDMhyECWTqyS5nkVy/rCS5HzMGTwF9JZPLUV8XoqR1lzPhmfzoga1aBgoIy2AfabYT87QQr
4wIE5IM1wSjJsKvarOte5EbfltXbxGKMCsY5BzUK7N2UrTqMI1WHGzvWKdmRMA91GKwnWzXkbGmy
OacOLnwr0kCgZjYu8rHQroSj49yzrHqH1pvXQKYp+9dFeD91lFNZR1el2v8wivm96dy6exQT3Pif
uKNjzLMJuxAPK1p+QYvdJTcw175GtRAiTEuF+D/Hat/rJJtIy++hePu8K5R45CFDYwaBJ6BLenpV
t+fX+3ozNoF+sbU0A0f16H4UTMCJqFZburtcPkopa0FWtw/lDcZz20Cas3V2tjzC0Bh6HvcMcd9s
s+rTHcS+DQq5qxqOt3wqhDM4arvPffm39sFtCWwt63vi+sMGB0kwG7mYC32XkazMzUEY9FTmSx12
ufCvM6LG0CV7YdZ1avM6jmRUmaV4Sb2XKBxKQP/wFIzO96Eux5U5Vfk4hI6Lpq7y/B8wJjDQTSf6
lJ+oQ91AvO+G0Ta0jpdSxCzn1wtLwICBJuYhR8l3G62VuVsoXg5cdGO3DrvfsZ7N6CiExksfyQBw
T8ldjM0aotndSJ0hTjio3124WrmF4WiuKQelZsy/DpU1EwiFOk6Cm0COn4dDHAVFvjdmjrai+6vB
O00mLYMojWlik+SgZuN8xKLuV7FIy4Pdi1W1ouKAhNUoBGFzQyPipK3SA4KNB7BLd8CEC4sPAtT0
eS9BgOQAMuTazsesRaNc/Mp9WKgc5MFx7Fw5/3bUk+DJ4/1DtHKsir0BPgho2fFR08d9DC5mDhEI
vBhKLtA4/vLIJaAPOLaJGM2D6BboX4CN8dEIzW2++68KUA0mKhGoDL0rxJG2bRqIUl7adD5NHXS3
UdHS8DfuPoGSJ7ERuUBMNWEIq4nRml3Ei6IXjaBHABYkgMtgxOASYVYnMS9Ag+T7H8O6TUxHAQsZ
iaIT8H6rJEOlxwyJt96u5XjzMmTC198UThlYeBpRF02zVn+egGQWp9OpfX3MffsminSMM3rpbfN9
tl0wC0EAs8JNE0h/vfhdZ297m8A8GbhQ04rHXXBqdruou0oZ578bMBA7UnC+k3Y4Wt6YXzV/ujQI
djiZWiFVWVVW4ePPqfxf2bv8c++uj3IhbiDlRi07QDaiZ9whTCjVJsCxO+uvwvfWqcBnh3lVRAsP
wi+AwtyUh4cQ8FYuoUeQBTJQ0QDHt8WnX/jgd/n30fQ/oJ05G3oc+WJ7kNC4CqHrFWhZaXmX4K33
fkSIecsQG2nqkx2TgPeklVSi8D1K/cUDki46gIVQdI1OdxzySJEirASuuHpe7ZntRuFZRCTzKqNJ
22KE+3aHZQXDaE6G82Ky5DP979qc0Dq59hF04+FMn2yegpMcQlf8VchiwrqE0L3Vs2XpW+uK8Eo5
+KQcYtjMHcJEHXcbWJG3vgtHTlUl5caNd6AJ2Ck8sDukd4PkFZKPcXQFBRugOD64tifx06PmUdSu
vQeJXX9Soj9kav5p2IMUKxnOaq4s0yk1J4q9jBljOX+UQeacM5DotBJ4BER+V6qQ3dMREH1KqDrx
JvavVQjo0kpZDKR/F9RYPgVvMZZNz04HYEibVQoPfBrZgr/TyRwRSRYEDwi2dO1A4oUteD0TSy7O
eRO0wQnUzjAXiCcddpqowPa1wgTPIV+8vqqgrJDf9anWJhqWcmxIM1/pdCrHdjLeKz9EVgmv/ehP
nEAbZocPcM6EWGoVsP0shYpL1Oyh2ElRS56otPZ7vBA/1pcdrycQmnGO9GpW4P5vkneaIOrIb936
WzGXH5eQNAzkHu/XXjHqu1JG9jKINIar+3NqMiOL4+4K0iH/TU6Ex6oNiS2ltGJ6bYaJSXABT2j7
gK3CymbhDjNnY1Z4rPyBndckx+S/5jL6nVqIOnQPnhlUrMpDCIRzZxT0AMFMBYyErUgZm6aqnfoH
q+j+KOFSmXmTe1Xj0O0Ibac1dwx0le4la8hYvGceQjXv+7UGFZ8KGBPkOmYEWwzGq6VcWj/43pFA
mP1LWg+WXSw5F01brb5xbbNr04mBA5CiRcSVYMW1iUwi2osRQ748ti/FoWbEEkcvt9jwTmlRhdjH
0Dhdx6em0XbPbzLTX3FMbt+nrztwczA58jSdGoHnJGMhdtYbngXrhSiFOJfya1faTGSigmwZdIHH
1mvFW6kRcStR/WrgRhqdiTGl4ARXRfh+k5Eey5Ham/FZFyWeGLTvABD1wxYTA6o6rJJ73DgjQ87D
KATF5Q1PNI3Wfy9++BqH/JmHycFkU/zwfX2VveV00RfdxtRkmONLPYk9wydZYgEZ/84pc0Zr4BqI
KRpfdnDkpLS8uSdzcaz9zl4fWDKQAkM4sRsCCvjwnFwasQIXNdm3aNe04FYS25PG8dCJkXznmhnR
b3DM3JaKatn88EPCD+jrLM+BwImMz6HUXYc3ZY8jWDHWBC8ajxZFe1/3jSJgC0JPxRGP2oeibtX/
Xx6b4Y4tc4AtEWrBCSsOfWXwyDa7QDs/c6iPvk5rmSNBpdA9G1z2j++tdx/nyz7/JroYP6XVglhw
PDUaEAl8Ki826G9OVvRhVjd4NUcYC6Q3rRQyKtS9nGt55uLic8q6W/POIzUR/P+oBIU/ebXN+VmZ
/ClH8GFDFWsLlU+Uj2LBHX7WTM/aCG0Dwjr13V7EALqibj3RQrf1+P3gO+4PvaQIw43mM6ni671y
iQbyC743IM+Al5jKgvu7QTgfF6ML/68lIFdLHNccCeuMNn+FRgc0L/R/MQgMqcV9RaKsL1J+q+EP
7Ilu0lv8tjpK0PF5XAh86rti+j9sqY99tbWZzh+Vy9TLn+TgJGg6d5JcSBKhFd6C5N66j4sllBrl
0d6eSuQlqp5dHVWmCs+2uO/NbAngOsaWVJyle3P4Mr7CSjVdLkRnkBMjTuvO3Sm6iV8F4mxM74p+
wo7hhKoIqwRywrVvMPoJYLxC18udP+U8i4caaGHc9NxtpkzNoWcpEdV/gEt8EbP5lY5CBTQVEKSF
t55VfwfMsbTtUNb8MhbefAnkJHTQr1wlLIkGbf574YVmImt93KYr7S011KGD8xWdjBqarbDOP8qB
KRBI2ZrW9Vqh559biNEBHnIr47q9dmlHhtSx6Dz1HQWakl1DrjYaK3P/FiefYV39Jp+atzhUdCGx
Ky2GVACJ+MInjGe5k57yR2K+36DlOz+MEyxyiYBa1efolquT98q4blNWRl1dqQFlxf9UKROJqQrj
YW4qc3tSIWnV38lKszx2+oFvNwmHbbfis7BhhEWqh5dDK9JyS/73ztpoupMbnnLfTeezWAZn6NJp
8HGRCB2ECHnkI8IUSL5v8MzRlf/s+o5k32jAbx8fz420Pgc3OZXPlxW4+JmdXg9xUXVJfCTLiuon
B3VXxUm+PZMnySXMfdSBqrQUT3CRRKaI4z2F8lAxdLzqOr8BBLERskGkpqOJTdCY1xghGKTHlq6h
AcY88dZPHfIWeG3/KtzmPtGqcsAN3eRFTHvdrTzZUO4nV+ODXgyfhsZT7sfm3iEEtzejEPMfFlut
IDmHxaJ/YgYxsuE9thOnVCy8B8bH5cB2WompH6AgCemE8ufQsxIrIKIQnrC1hw58Vrj0JhmBYJcp
/rD1ZM20+KwQy2rcnjPLibpHJ6AGDiRrqEnQr0lDEvPUkGsBGcP9js4l7oamixu+STdrgH/anMhG
Rbh19L98SjLiXGUPyEdYRYTkoBl7nMCb72RBAT8y/xqn2JwGhCGBK+REj96dmbfg18nUSKptIJvf
XjqnfhHCibr1lb7/pgLgoGSc7vNX2CW+85TtK05UZ4cu9Kir0QR3qH/hRL+HMz4T/obzG4w4QTrB
PQ1MAXnQqnBunwExdfnF9SCyT+UsKRdaio6R33NRTN9/BvDjyMprmSGoq8G0kjJeIeQFGyRrlzHy
kD0IfpBFINHFK87QHWs5HV1aqsl9kNm2KaxpDBDGBNRTnJEZfrC4FItf0N2RV6pr7/GWiCQ5ddWP
uPHaKe06iHVF//41lFPvJAMMsk3gzIDYnNbzxw/kIN+UPO2KGHzLiOGeNlmWYhmNV7JYkdQLYIW/
PBxVRJvHT09eCJQGUblUQ1k+IgghbvsaUO0WmUzisXvpVev0SC3TWsgm6/lTuOnmeyEBiM0oJD7l
Q1WIE+DyxnsASCO11bCBDI1Px/7j7TEE+jQ7xYKDDsb8J0VVgWmRkJ9+twEzUrOXYJ7E2x+2ubBz
2BJ8pwKBKEt5mWw9KmC8VLk0E9Rlzlm9AQefd0ZLr/wlPiV1BU2Yni+hA5hXDvXDYK1AylxRzvDU
h/ccbPfHZX2kS/zmwTJGDz5iqrDRWIQlgTVK/YjovWd1oRfpk95yWqyZV1JbJ2bj/L5TLL6WmL7a
kpDLjqazKOCb424ZT18L869rRyP0PaVLZE4/Y20bx0xduydjHvTcLfMB289W3W3lEgqHZj9exIL7
Dig1j6kI99+HB0nidJF4iXlvpKZQVug7fT4OfLNtM3plKNhm2SImXtmQ1MV+0+nG9aoesf2TbqSc
o11HKIW9NUO4fXzA47YtR9Bur8gej2xf4YhMuYU7PnZ/hDizoFVVI9gKb2YXpAsKJnvfjfMPtCAy
dfv8X2iZyQdcRuwWgXdS7ztwVuFVkR7ocL80K5s+uu507r6MiHjUKh6+xKqaktVzOZlPrjwzN9Uc
ENvoQosLx/Oln8WIL0+d071vdlNfKNsEOB3nh33ReiWPC4PxvMg43ldIbrLjNAOxk6/mVtTUkuC3
UczoKFDM01wBfNTQ3X3rEG37Vij2PukBP2mYR4dS1+scIUmp/dcucA03zkxGD2JO/ayzX5qZfc70
3mujm+Mhk+1Y+Qaq0Di2kSnR2t5dxjc0efoUGQgby53bMkDYwaNOURvfJJUe6qhbOF5wQBbq6yL6
nNNSLJZEmTmwmSI8NRfo5xgzs5nypseU8YQczPZ9aj2DY6oRfBa5miaNJRgugfbTvWIVWb0r67Ec
tvCi61WVxPcbguHpawIUcsQufRQe7aQEwi0WNEb6Ez61NtTQRoJKrKrkUw5WJZpREiwh1Mh+4/cc
tnLhH047mcfJQ2m+YyBVyO/RAR/nD3R7Y7L0dmkqLGcsn99c4WIp6y40djQxa3TKZ9hRZF7d4rV2
34E+w3AtrGhtOl4b2OVT+0B5t52exKgYLM+vt2S1g09TxPhM4LCneFy8sYGuiNNUBNKHCmDheN1Y
Bz/gjyzWMHpea83JNomC0aYk8H7yYKf7E8kBva8oyhnis3a6qlP691ujS69Sop0DEKhotnf1KVvV
T39gVI7f5VAtfnZWsp7jyBvxbg0jDBUFCictM+hJndbFw96MJi5kH22YM2Kj7GAmbl/RR2K0kSED
gmjJbvz1HF1S1bb/ismkQXZ15gl6VpI6kX30OmsnsaClXh9eGZunz3bz1N2mko0T3sFd3QPjx3eC
mkJl7DXCGu2sdDp6nHMTXcruirV5WkfVkrty8q42Iea6LtWcG20bOB6xEZmFCY8SMJ7OQLGcuxTw
WI4Eq9B4z2Y4iJuGQ2SMlnrAuftwkQXrlyZM+70KR9yyEFtYMAvBe8mto2VgwohWPJHm6gTTQlpT
aDLuMLcjnBVrFHCFur+cqefhnj4ozswd8gRZAjzTSYoGDJzyIHAN+1CTgQGNy3vhDZLsPy4UVMqK
Uh7Gec1NWfc5cl0A4ku8uwypWq1zeINL/gBVD6wBYPRGtDw62aOpunFiH26Ysot6KXfMuH+TovsD
bkGIXaxTnEaMvoVZlGrdyOit4P1zealujwMlwo0lZRkOATxgVCIGPXz6CbFyIn+YzUewk9EoHbZB
/JJ+ezMPMGkwPrnMEy/TlGGig1kobZEmu8tNLyOb5elqEOPg760JJAvo3rJ4UP3AMmzrck2+PezX
dLgKbMlBTbaviCdRNPmfoIlL3I3sLtD7sGIRTYF1eJJhm/mNkst6/XTbzCxe3HE42IVOh1Oh5/um
T8fmvxPCqWY9PpySGmmBtQc2EkYeu7cLSudH7JA75/sEQYT0XM76x0+wnwi+hCS3ZRQrZOKzWnzO
FYka1r7ATTFqp/r/Bl4rY5I5GUGfRu7oa1C7FiUJaNhk+paEFYmRtwXNxx+gZKLAlnsyrInoBQAd
lGVAtBhrdiitupg+WBQHNO0v+TIWJPPjDQ6NSXw1odOkl5x/zISFdWd842GtCO7uuXIeUVg+V51L
4bKtAOQ29ik02h/hJxGZMYTItik/Fzhx3951nu1xbYU+yAyLxoxyI5RqKOwOvhCRV7ceRE/zSXyj
LPYAzBTVfSzAaSyB7oKLdDsYxvPPQGG/+sfxOHtAABpkqo9nWLYZZ2FytgrutOZKJgHLY2toT82v
TfrwV2SknGVHS8Yc0M6GvxV/EoYLcnyceuqApyMhlsQL87F5/KumsVYAPkcor6/XUa1BhPCTtDiD
/9xPFImpXml8oHcWd0dJOfTXQnoyI4c4bwCMoJP7J6Fm7WZyZwyP3snIqlyOVsdylj8EPAfplEMD
XrY5LWFuyKC2lVQz7gLe2c2xzVAJbULSagmnGAJR3D+HpcvJ/C9PYPhhwHF32JaXVqpsW4Ya9BBb
cHbLwXqJ3/goDicZ94JggOI9A6MCp2WHn6uiMGS7r1A/VJP0U/mwyFw0eMGZ005RanAtVZ50HmjS
3G7ZtmyFzOChvgtgm624vrAX4SVzeeSFDIByfkdSV/9GvMAJ/E/uyOj8fgSXzJsFua0Q2T01jyja
jz1UMd8187OvaIQxFiXSjUnNsRGN1qkCiZW3tYCM7/v3VHd0Vf2LwUSM6xSMPdp+sU3R3uJN12+e
HkZU5Uz3p4OdYV0ImgOgOP2JfiTXWiKYvGU9+mZ3bi+SqYy5saCvLak8je13i8VeYKkfPECMSHQi
dBa465A4n8+jNA5tjN7gYkeyIAhkhIuGz9HnNXNiboBQz0ojRaLyOhZ4vRjLoSZOOXAYhGOJhkxi
sdlaZTyh3agHxS6uIeYs33F5BaIQQBT6LYi2L87huaZlPVOTYhh2uERwcm3qB6pkrw4m+uJbQlTS
lkTLzAzbxqf2TJ0dGv8EtD1uuxu7r9MzpgfjsMECh2qgeOYVKj0+wUyrbV/R8+kEY44L5m+vn1rT
qw1d39EEhE886EGet+9PjwEKUi7G/oEMMm2jFid75RcQBW2KCC3HRB3uJwdYokd7fDJfAAxIzmCA
0ePPWL8Dcy600u3OaoqBo27ABIhBUKGXiUjvKCPSbVP45WlaGD8W4GdUoNnjnosLkJ5EyuY7C/7s
DZVkeiNR/YCo4kJ4LO9ZedIgOG1HkdwUFsBfAD7Jahp88pltayDdu0W3GsR9hid0tRyLwniORMq8
UEj9glQ18C3OgcThB68+jKLntSXD1F7RZrxJ8JbPS16LDDS7t04QTwzq4/OFPV4D9RYrTCBqsUcl
JuLKMcurOSScC2xmi1r5+6pjV7EqWtlJTEuHepZFHjGcOnCFISgX+tzs/d08qibME4BUyfyTR7h7
pwiCKwYuIX/dEMbujhL8USScbQXKo7aUN1o28146wmepfiNGAl3RjQxFwucZAkEajYL6nmHzpbio
1wctgfcuwgWg8nzj99edVpBj0UfRYMo4/SN2R5S9mz9YPxhgDDnn3cgmHRuZMf6bvAUVnLLiFOII
eQVxToeC1fhE6UZk9Ix5fSDGHJoLx9uxkVVnvVVrmuzSsPTPPlx9yNG5IRO3mFxBiUmqOrWIwrKH
9l5U4+lT7tsNa1WjSRdOkfJy7v2W5h+GitQK4yK4yM1IOpDOPkntG+1f54Uu8s8CxYZv8D4F+nfS
eKpvxQ3qML/d6AOYgIM9PEsnFeLbrP8tekoAyVWo11xHZSq0V8udMRAByi9GDaiXzKTPlqc6o4Pj
Efj/UBMoZAQqL63PtknShUMgwz0NIA/rFGI4oKscmSGxknrI3UNFZapSb6GSqbtqps2qManJaDnU
wLJi4/U/YD400MPR02jtT9JYEPsUSGCnYXU8ascf52Bk11zSbEVZJAK8qfmA4gcoMbb3K/nmnj9F
qutdImUejcgIaXtg71GdoiLfdJFM8ivrn+GZrA6iC+gh/pHNFHWEhSpiBe2PGmCaoG9Kk1e80Asi
O7JBbq83XJc36svrWC96h1jJjA+rZqdOB9cEQvcFWLSfhue2NowK+K82Rkxzt8kFth6spL/x6vsQ
6z/ITgeVxCwvwpdgnK/vxrsY+ZyxQ6DgZ8dF56xtEg6dS1Kwf91oQrqQlF8h83txcfn0MUXwPz41
dOZEg2PQ1S5KIelrqfENsC4Pu2J9bdnFoUAFfHL/g3iC4AXqP59vRXW0xnaVhTZ7hEL9K0Lo6mNn
sHPjh1eI76IwRybr1g8aUN1vxgxuSr/GfxyaoBUiNw19b/V0yBMdHwFop/+ADlQsyBEL9yQsc5p/
xYMrGznk2pQ9lW+aDllX4B/kQV0B6zwqFGBCX+bZf0fegP9/AH9E+mSMmWydAYO3oBs2Ri4Sh1zj
vuyAGUol6/4N2YusSjY4Fig3qqlE46jY2udpc7EQ6sK2vM0aeMtXzKQQcFto3BpbNecMv6MN+FXc
q3Sdt1h8K1NFhjlCsCGHdxPm4uVcXa5MmihPDypKNS9y+d+OfFm+f3Dz7fjCAwQubc5RXAbOgF+E
IvEfuVbjM7TdgpyjJVl5XB73NPIpdPnqFY5NtsNDEzTSRPfTARp19L7LSnvz/aXLJr520Dvx+oay
lKWqXzobQkrf2KGzKkuXfIAuYha6hEvcEQ9yImvdoYmIy5glAZNtBckyJviCrLuE0wDQaiVvQ3ZA
NsKqTlIxZDkoyoGdtsLZA/DrizImz4nM37Pp8HQMY2n/mjF+r5oCyAp5+MBiZdOZ16CvWmS6xklM
njs5PY2u3uDPfKgXY+eWhLERL04WLyLF/Svi+LDD2/OInEQnB99EcGsiZBZtqlScIO9CeqeLo8zY
J4RMXE7k0n6/9zqkOc5160MaYocAv8Ep2u5rgzcwYXF0IZTcmakq6fG9nG6bZ+Y7EOlShbJLk+RA
3HXhuJrnlcml3xmZNNyneH8qQulQ3VER8z7CM82x9TxcuFo57XdeMjAZKxBcCmOZVVfs+yWTDzfU
/7hoJW9rbQKT8KYs6GiUMM3TZhcj7ZE2NPwRePuM0mktk0loOQhYoIN13hYhzBuIefi8kvsRGwvE
NiB/06GVRtwVYGZnYXYJsQpxweZhJNI1NoJydrKx5ZSWBFffSaNrIqDJBR5raR9aQDRzHymmV7t8
qo73sU0hOLAAqTgg6LNoPv6NC/OTgxJpYodA9CkRJox3h0XToYMiD7/U7sCPXSjIzUWSMVNMiIto
BtnRfbO0Xv1g6ENc/aWnrHtGGZR08wRhWAqa94dlhVhpD5nFZOndshWS0C1IySjSLHtzLxXgRknJ
lhBZLRvHalu2WudXZKjzIuMD5LCELByFkzjxWfXH1I1QCOCxBYLfRTcY9o4MnamAioEdNeA7Vb2Q
SlyOtgoaCUHc0VlDsVjf3Ft+ILEoDAP1bD29TSTY5yIFjhZcP5iT0i0ss0nSIlfidNmruJuNnUM/
E9sdcN/c/Kcg85rfAiLXLba2OtlV2l8z4CiCTskgR5M/xUFXMC28sQUZYXGjQb8D6nSwRxSPWnDY
HErOHDVeJr54JXSt4zkbpm2GzqnL0HIear0jcNqtxzcnmQPeJAWieSeJK4exMqa220Ajn7LOjl1W
UMLdDtNKIiW7HW4oA/gvi2917E7p4nLN4GuPrexNNMMsj2kVKWFrwV9hCujDQ7PCVasSjxW9hXcq
v14fjfgpMizzotmcWePB5k6OOXaoOi1dM66g5CjgZCX1pyADW73EXtGZr8y7a7jjjr2hNuXHCo1T
Op5PSPutZ6BKunQRi0F8KI/clhctrs6HiqmL9zdtgJfYgtpZ33vPJpluz7/RNVmOrSxQanRd5Qlq
DuX1tO0FBOpK61ngxhmOIaiJZZhaAFYFs9KfGn5t1eFQ2D8AzKtr9elIQGGJbFCK3/8C/RaDmj1X
oocC/HMuswpUSM/5ipH4SZvg5g3FjxbgLRE8kIITmE4QIOMAtvJCVRShEQK4Ur/2fxLWpDdQqZrS
CkHnjN+CJinINnbOUm8rL+Sy7svvGsUa3EOqSqFNkjE6s+0lgg+1chaqTNN28sIa/b0OIRRNXhgs
MvxHfd61QhRxBzaQ6QK6xBqZqbdDxF7og8zFYlHgkfg+7sbSL4N9EQxzwl60Vu6iKIUNm68EKVbW
vMHNjzdu09g36JwRzu1BBMHWsf0YG8Y0MX3Jxyp3T5rq3H9T1qMG+PuC+Yuia++SUq7WM0xEu/5G
DdlXhxWIe60Yz+ynyq9fifShdFS/sDVdv6gQ+6src//NopYO70JgXo10ZkalOFSWPfPsUiINa580
1F0VeVaoIS4Lg90/unx73I/w8nKVNtR+t67xV1uTkGO6QOspGVOTZm3Tt3IV0flPjq4WJPWkRVDg
MXHskk6leP8DQOfp5SZ3GW5EXOSUDPi3Sm9vzwnbs0bwtyl75Isc9wdUS05ansZ4WRu74A/LfKzZ
dUJX4PNfQsaA1i+j8Px4HwpHavuRJmLMvsULJ/j+cODn0vZk3COETe+Ot0b0Vwq+vQZYsmK0/eBv
u64/p5V8H4ZG9KHrYgCU3NhbNV6QfxHq0qJPrLk+IUCHud865A9Vz2Ugu8j83z1NwH0QpRxqZ2kO
wYYIhz4aVKHmsoNoqyyeYHurBBlkGp+tmHn4PjFtt1RXSSVl9FiyLOOfV788U9zGEEOn/mgjSjLL
6EIAbYvu4MHHMKhfSh8sf6ZrIraSDZLMpFn16giLojJv2Yf/fqTtFCckjt8BUKR5ntt/kH5FAerb
kYI2GqYy7zoZd6dh5Sr6FpRByCJp9Dec5htktiUhjB1GhpdW7zmtOFXOYt2U4hreAZaoBsgJLWGT
MdgNe2jg3CHqasOxXbxu0mLVgkBRiwTeRtJkPBKP+PRXdhzk2BsEjEtH4A9ogju36YEuK1PFeTAJ
MnwRR2CD9vejc3GkJWFn2HRAHS5jCRmA2gnHDeVs/XBuFYIUC9PtOOkaQOAoQ1bM8UrenZvjpiQd
RGpJCieXPxuo3sEe2Ln0SOdtxeKDQn7VxmYbyVFECHaRzDOIzKa8dcj3VFlP7lir0RgW5gULA01g
BAkkkqOfJ0OjXDlhoq7wadcrvjeLd25NMJZ9LjPjilnnNPnOXVijlGuSGZu+7y5ryfCqv7dtqAww
KvmC056lyeXHnOFkvNoVJVpp772EfseINpxZ245Jl+jgz3234XUNnxXY+yFHv8K316qryo79v0Mc
jF0nhVD5BzYYH2kkGMoDz9jWlA0YgZe8PZhYYpqpdybK673TTO/vfvNbw66aKDDbEAK4YextsbbN
BwdRncluLYAUfH5q+L4sz3cRSjonhrOWMpFwGUReWC0DNRiHZxsFM8gUfkkKMp9MUkCOrNhI2zGh
rOMBCF5m2zrmJoSGSa6waWsTPNe93bpGvddyaVOpsvDTJdUCvvRB06DnJiMOrz63Hc7uYiJ/uQuy
MJY4W3oUq/Gfmc52li/kpFO/sYuEC6jfGBrBamt6Tn6wYRNAmY02hAs5bwln37MEwGwzJsdn7Z/R
nRKYzuKLS8Ca21Ss1awdlWQDwKKhVP+ZmsGNmF7fVqdILQV7IxmNaKtWP4mbE9jbSaL17gZcOJ40
IPtZNvVho9DCAsbkYa/bVv23VAd1cvzv9hcx1YDHFLpNcrNr4paeVynSTfFVCQAM36ap+4SeAL6V
erHtPBj/i9fVPE6HA19L/mrocA1bBOcvLwkn7pFt/0jCQpmt0aDCh6YY8sv0s7+iGChjScAjI6iL
jK0YDsQo+uXQaj+8ozYWLkDgbgVn+PyXAuYvYDNARTAFpIT1t3A7A5bR3ENi7Z/qz02b30n8KxMV
PzMYODziLiK0ZLoFxmH4Iq6frzjhHaN4ZEjzBw9Nz8p1yRvoTnZYGM36xivNWjK4+cik7mUB1QET
/h435s+le0YgpA+YWwU2s3cODS233uCH2kF4Rfu5IbduOiAPxwcPKF3us5RKFUgq9yMct4p4xxFH
H37pjIXQGqpLdVimUw0eG7fCrqlp25Qi7VBwqwJliO3vMbMX5h/FQH8PZ1VWHHxKPuM6GWYVHdUR
ulJVSxALy3yke13DveTJRJ+P9MlUBdNWv+qMC7S5LSfuqzIzEYqe1viiLBspEK0nTQFgqH0Q5Fb6
mW03+0sqOuBMj2cEEKogjrKWeii6+Os4PaaqV5nBa/08HQneoeIvwGmljQzfYEVt1drwtbIim4qT
+zNqtXJggyUc8l3UNcvOmrUZpDjWcKmM1EdujUfr4Nvx/C53l09vnJpw4YdfL6o5I/Pz32wp5Egi
CeiVwRGMkPGDzv3daQXkWqsQ6m7yaDBMK7jtv05d0UdP+jE55uSURJZLMyTSepXp0LYQdNPkOLdl
URL4ijwdBGmaZkrc1WWcKrrnxR969ihBFVfPMKPL9ShjmRKttu0+0lksd0+gXjB5kmeCms7icd0A
8vRkq8/Lx8aLV0yDTThKjLQy6mQSIaPM3b4tdvjdvOPOXYNnxuLPVMoFku//gT3OVSrhK2392wor
0iKBOMqGmpI4DByrLagag7L3QBcbi3dLccGbJIdiub/qlk/6WSMSLynMP/xFlXwKQZIiKt/cMxJy
Najij6c3G85E5RHOZN/E4md2dLredUrf7lNZ+dQiLNR9DRWqpnxMomEFbn5NU+uosZPiDy0YRh0Z
lx9ybmKfFvPsMCWbiWdNFD9yEdwOcqAABfgjmbzQ0cyl9Wk439VaE+Etg7f6KZ1F83RbsQQP+/58
w4Pdcc+jj8gl+2u//b9944Ria2S8haoh79MnRvSwZQZv/UfvrN7NbCYZmAg6r4JkyvI4hZvdu66m
ktEYc3wnWeF9m11cFjff8WLMWq6X7Ocl1QaSsX1n2zF5sx+i+ozZS4cAFmZEdLZeXQYErBHMj1d8
oM5Sojc0OhcZdUir/g0R/CkhPPQYkluMNQymSFOGCRTdPUrcguv5ypKyLWllGupggIAgfpQXaREK
DmB/R2W5cNZCP5H7OLSGXuYrhUcG/3MFHp5RB5VvonKvhEdUykmsOinokkOF+k16nZ3oj8LnD2gf
647vHcVDovcNHdHGTj1uKHTRjQHtfk6yfzKDhrnYMX748eQxjdAL5utBR2aM9mpChZ9wABguipzI
Nf7HOxGYAxnqnxzGoIpZUe1/wUs16SfjxuahMCOQym3xKfTj5uDEWn7g//PLt0g6JeRb/VyLXN0R
Ke7A2scuCULUJIbx2aCzMI2F8gNQLQloCWNLtnbAwvWd45s3e3yxefTv6tPBQltuxnCYv+k+S8mT
g4EEZRgaTxMtVnriGpp4W3BKE6hk9Tojxibfcm2I9AuFxpzjYFL1dhMWTcuVYuRgNY7m8RW6sFX1
1UZp6TAXDjHHry7exOxrowctTArosqtbzKj8nFoaklQowpF8qzh5fThQvqIS0IvxDWsf5ps4kIFR
Qy4GdZPGVWBtmyJMfu0Vk5g5Vg+AV5PzW7vuvbv3I36XwLONhZR5prtOCegGLKgcIN7OUBobTTvQ
5VdT5/0aLmN3fIMjmQiaTbkwPKaqOufH1o8X4o2zcRBlVPBoA+Pc4/iUP5Sn+iDHcChUsaESO7I7
Ypc74LEJzG7AQod7rKl82IB177TYyKvnZptQ8J2XBISNjEM4Rw8J3dEq3XTmlKxu3OS7b2WUg/Xw
HukL7ECPopiXToShcONf82kft46Ik1+uKR9p9E8mcbRxeV2zQ0QdEFC4UWwBJfOwww02ECbvrKfT
i0eIubh91YcTyJh8cbQ0pzX1cy5uL1LcQ75RNtUhyDmMndcqtujU6WIsfN0ti/ExQvoTH+r4um2E
rdjc1aQdaYZDOaSy2bdfcCSZlNMx4l27R5Rf5Gw3lxrlr4kRRojbAfGJoC/OO5e3oFZAOerA97KE
Eq9wc+RBjfZJKhrABe271FbKYJWvwLXHrub7GHjLbAhGK4q0n8VhXu2j2aumXMcpO7//wcMRxKPJ
yMkkzostVq0fWWc9bxp7PHYfLBtsj14b5I27XH/IjiMCRP34KchpqGC2Ga+2csXS8to3ij4tGhk8
ts7jKlx6jX3EvRk9GsF5S1sLGygdqNAU1/uXbV6HNzhwLGgPowPtQUE2vC5f4JT8eBKMeGTVu8xF
lEDcp8eJujBlC/5BouYQwlT8Ck73Xs69WDJx9QWt+qgapUx4nzHRQ7fTykQvPoQHmDR/J9ah5uSL
/f/tRBOQT7wnwYWAcLqSC9SxjrrDE9DqkG1IByKW9Po/HlAjJpWZN4AvsJE2juXFZXFUAJ/J+8R6
muI4OPLksbUVn4WT6rBw5EVcmDNGFxMOiT/HZL8pjsFrNN/f241c+L7/hG/HBfp5juWjCI18uBu1
75pfWmZh4zG5RGihXc0+k9xJJ0vWdsLWRuXCy/lHNrYsuYDqOSeuPTcX8VyRMX9EFtdUJzpkf+CH
gpxXH5zGWt2dguU7oxtCwhVlBZGgpzMv8WYS+rRRXkdo5eUMYTkqJ44Lv0OgpXRLaGDJxO6yXcpu
346OynBYPcqsyyOOIu6SgtMqfgc1IF6STV/fz8TFA42rfpW1bM46LoP4fPusUR4cVUbv7tI2WFrd
IkQiLsn8EhYkTCoOUHuedLNDGd1WxyX5iPDhL0HKT7rt1bkcQkpGVHklP94+xV5eZcst0t59t1ph
ossZSM7WaVP0Yx/k55fvCO0zz6HMMgY/6zl83Hwzsg2G1vOpUJ1yt3ZycgvLLqnCJOWRPNiN/ABc
4U8AxsK8R9zWyoIj1O2lLuWGVZsaqpcBsv/P7SuetwxwyGWuvLRUE46R5t8ckmpWYjDCjjauedoN
HKbU4LlOVjEvD9vbuZN27DhoOJbJZvSk4dsHG3j5kCJAsSE1tzPwMZRPUI0otKEigLsNs80ySqaI
hhQdtYZ8kXDVyDtcxZCYMTZv/jQlFAJIUHgqNOizd+j5CtviH3t9F1ZM5beF4VA2ocF4gRpZz+he
sc7zpRfjs+f0zCc/hNsSXSGBmvrH1uQ76RWZU3n1bSYnU9CmBN2hHSM0ZiGHgpWjACkHlavI/bfj
HnqxNe1ymq/UKpEMqDAJRxyVYsYfz3FsBZFjVPj7V6YTOClivsvGVJddNvUKfuyqAuOyTvUNr9pA
DVhz7YGWDErjL0GKFBb0/gF1zTbvAnvAT2tY2uSus/jBLJuK4xpaaLsM9qjoVnCdV4mSBOHlkQXV
fsuHi6r2/IDwF0FXHegTXfmohinWMHvpOSVc5Hqof4bv2liQZPC1GdwTxWzl2g8bevTYzTmi/Uy/
fc4uaEXUyGfP6fZEUJprPNw5rSOSqJHpgoBo58oFmmxxwctLS/RS85Tc7r4bQl60unBexsvZzHJJ
NdgqrC35KvyRyAiD/AT3Qp7vVql8L0iq+UzbOrFRQiU0EvLHrNdvlfyBW/VRlyx1tzDJGASEg3su
69BVrNg/2HZmD6gIDZVZb6mK6q+S7T+Pi1KpOwTw8BPgeFdRkcVyNXVzMqiVehbuN6kUeHm7DYpL
dYCPpjWTWqhNR8wFNVa8bEEG/UBmJoJtXcwExDdAQu1lT6p56HPyAJ8zlnfFRdtom0e9YiWogO62
LyUC6aANL/Te3L0bZaCVX5OdSqKHMGzGbD9zYn6xOy9OzJjgEsDO82FLDMIYbS7hhVj4o3kdK9FY
/eZ3MCwfrwgfDieBj9L405X6k/BRR+Ei/frzPdSqWjisTQoWxDurqvnbHCcBJJ2s5yTUXQkZ/peS
lQK/i+kXWbroh255dDkcv2vMhzFzkhko2ES3bLsBsDuCEe7i4lK2H/fUFWJZoueV8Ix0MQd+lRIv
z66rP9+LJBa0dQ7ehAjWp494YNgbQhJBysxISroHcLygZKVZZTj0MEJ5OO3FcqJWVBJhDnPYkALa
aIPrfBaQMNXGoVcuqe45gBp/C8xpbeNljXJakLakpJpcGi7DR2GNW+Zq/1+Y0rdm1laOYFkiahH+
Amos/thAtCPIgb3G5E/IZMCupjLFDWiYs8pWmyMBCbIOikRKKaO03xkMCU5jKicw7Y+3pcJ5rcdX
skXD9u4jyUM1nptBePDdBVXVkRQxH1zh/+ZGoqgl2ukyL9ONP9X3GSX9nLs9e0oFVYS942phkCnV
WKfAGTc4/YFjESjjTYAiLyxrl54ZxSZWV4r8/q/2tlT1EZZfINmsHl0vjR/hiIpwRcQ5E+nPG/zt
Xyjg8+cVe0NQn3f+5TzRowhOLP3eISGTCJxTXbibU14iIyMlIB63s7iRoM7mPI+dXxRAIL2f9xF/
jvy/3AzLxBClAUB+2H7wBOqBNA15d3wH0No4/vbOgpXu4Q7BoFGgXJJ3Qj1tfcBepjjQpQmbklLI
gY7B9jiKSLhLPfBKh8xnZZkFS9JP+1s3nwQP+YVwWMht0ocAOhxJheSxnvBRfoUQ+Fl5vzwUr7MQ
J1k1WNY/5Fip952vNRqb4cRHci3hGTbeeoK9KF9ROg0jjPv2KdxG7K53RYkjSE9HN03ZS/80muQZ
sNfHg1oYXFElOvZz4gL2UKaHcMKygo0r481en6plFEAwwsz4pyuSE8yjboFaz0JnPLsqFKUNiU85
Cqpy6Y6EyX2oMVHjBtnGfbn7xu5N9aghF9siFgGZOYXVngkALOLyd/AmekxH6bcA/uhzzijMcrEm
uINDxLLPd4ILQ9QFoFC5tF8YxCguIhd8MBP0eZKDNXwsdzN00GynVlElIsGFwSsA5c9SG4fy656x
tnPFfYZRAcLw6r2WjeZK915HS+uFSoGiDCDGBbrp/kfHHsZSuVRGAPsiPN5v1RfhlrZPfVtBO4Qq
MLHQu7hdUvf/BZ+WVAhANi6YjDV3fNSOj2/QT1iIPG+xHbLYR54OEMipc6mqiJ2ctVBavGOfFmAZ
cE6dlNh5rMH2AHCXH1hTNwI18oyDOirpsdPIxk4Pp7t5hsrV/7p4eEznfg1WG92D9ZSAY7HDHjCo
Qk02rlDgB/Xnv4kfE99B5m14Icx/WjXARC/fV6EYczqQNGz9SHUC+vVzQxjusP6sUyj+dzUdQHy6
dCiroSaPSla5TuQEiyJxQ0CdpbZsNDDD3TEhoMTZRz872LQKcKAHkVzClQpEmKeHXS3rCudGJ+Df
l6VU6c9SN+8dBlw8uFP+Rn3LoH7o9d1kgqUU1wxBmFNl8OUV16kmKqveHRMLjs4OpNue0DHAAm2Y
bciNB/iTkngAY2oqD5dgHgXv3Mw3epBa7dqrGliglVVeTHf8VhFzZrUYNADyhrG65xEMhe5j6IpL
BliSJQL6APEWzB+4dGQGM+NL4gE8oq/ZJSRAtOQgH5ge0Nr1747nSu398rZ4nN5vb3eYxrKfhNln
nuk3itE2qoBL8kBjOc/HosvizFoBH5/e0J3WaWxZUGe/mR4SoI4cqh2f038ywXIo2i3Dgq2B0nCe
xrZPMPt31zdm68O0mejHVrDeTkoZQp5LxExtIatU+TSEcpzFP/elJLFfeDVjf9noBmpbSAhV5LE2
kKmYXQyYpSo+AjvrlTT+CvTXn4/DHmeJ0ZC9NC7NBAg1LDfpicV6QbqNMXlnnXdrWnXmWtSDV4ug
woI/wA91D8MjNBWBOLfICXrvCUL4JxHidFpZ9R92hh2UgOp1qx0LX5PBI29XeLaYtrnAF+B2120q
RG3KsF4/svKVs7IXsLymxC7R16TrWKcHI5ItIcrxDw7zGTke+kN3a6oOG352cErrBnvnBOsHzcG4
DhstLfZkvyRRtdN2JKDiWrQlQb3LQLbZMupHna4QVvcFRUQrvyLzU82Jm4i1OSJOT67P14BXHzzH
TuaJO5cEx15qeqL3vZPWCG6iepZytouwP7Hh2vn/tHnlPSPK7Owcw0XdfkbOQZ4FAa+4M8AJ8RS0
isp3FdTUc+XdJPAex0d6azYamCO07OgFs8oTmZWRTcR865BfcrygTI+PFEZ1Vn/h9fbB1MXL/Lxn
WPXLiNJYJVFozB3CCoMPDhKryDY7oXbU14+iF8s/Fhg82WOVuMT1oJNwLM7KVvswN22zb4mtfvMO
4e2DkrofBQUxsvysz9NK75GoomXgwkH07cz/UszjcwaYvPqeV9w1/wV8O9ocNI/Ly8D7xDxPsXTE
cHGbMDdy9GsBhMOoBv43JvnWzIvqcOMgCMJ0wsaCfUUB3bWrt08OsGEr7ezuG+SOBYsL+nOJvon9
HL43CyQ9LK/t7BtXsDNW298p7+2O1E/ZcLDpux2GPxl0lEGKCodf+T0STNd3lhUcIwFHY5ywwpI4
vQ+nOX2UEkyS59EmI9juf3AwftHKtDzCDssUNQRNMTSaViEr5r7nBbw9CP69fPmme3CNlRwPCtoq
lqhpGHbCNl3kND6f1QRx3vSTL1cxRHGQ77I46w3b9rmMxw0fVJ/YuProlj5ooe0dVRPz4zctFJOq
YwtocEsXHqosMUVfzPLZDCz8ufkCQSqcHzEI577gG5KSonWkWyff4rq3JpZKFJGm55J4YcxUiSzA
AXPrQc2MJVBqXI2EZFfe28Ba/V5dtqG+17eJikXbMqgm4Illq9mJpnz98Z/kvUIDxpvzhKDAKphB
Zgme8bUITD6rXX/Suh1YJL4aj+i3ZOkk12rp2mwHBDdJqBRn0WAiYL8+gUTDWwFVn3U93yzU6NJZ
gkdobS78SzkJ6pvOYHmhdc/NFxXF/KS6CqkAKbQ3FTBPgHHN30xCjd7t/nvgUw9Wwn8zrEXrVEXc
VfULGCpiW3ytDrIlOLlzQ033PLRxU9JE62xJu6WoZcJKatcVxQFSEnrAjJjnipg4nH2ma6oDxCRd
hxxndEZhzuNbd/CamVNuK8D8qFkkKHreYQYBhFhn2r7kB7cVEiJ/WvWuH0MY25XzcJir5irtQozE
T0bJ6qPGe1YbNeFQtSTmC7mMo1DTzJwO8wVN5zWbpXw8wSmuI44D4oPGUeLrtDDwdvmpGtaFyZUH
UmAijihiZzGkDxrjLYt7E8lHDlQHwNocfRJbRJI6e+BzKSAt8mDVx/0bgdwiOqL0hjunMCqbI7qD
IvKoe2F4/uOdZGH3rBUTV0I+ney6lM6aY0ATgr8wUXePkxyhS2YklLXep3mY1BKtrVkn7lZs35e2
ypBtP12gE3vtoCzWkuRjMRkg3ZHLzcIHDmjrfaM03S/jmcuBrGONJNtE8yxohncKG9i3EPrMcILJ
b71Chd1hRv2eyJKuvKUfvOA1puASqWfbUiNcZdFgw8/3nD8ZAOQC+M42TQolKbkgLciUUjab980a
IUwa5n9UI07uQx3bTPuY/yzvfOmJKjAbJChJR7IyyqzNT2JYoFMciO7l4peaszXMBNhZfw7ZxQ4T
9hYobvzv5tEcwlUUaI50Zll0B67fNY2j8T4c90UjEMnb7Ned2Atxca/xaY7WqqJJ9OKFmzifyFHK
vAiYPSkOVCIbM/j8S4nAhlkK4sZJ3Tc3vz2Tyi7QX3842N0dSeuLx4lrSBcHOvgJw278CMXD62Ob
6fddUEiBqoFE1r2qIYSTn4pA3UiEsuf0oYFUwREExK7NiZ4Rb7oN0wBQCL4mRFyx0yjM3gPPkJ33
5113pm0pV3kkr9Rf3V+Xus4qNYC8yjZGytKkBxjZNOKpJJAOsZmINYz9W/TgKf/SHaTSJ3cpk/ip
wHMq11e79FlN4WRX8vJZxnvo75bSzzrIYXaQuklAXAXq67wGYs6lsS5NX1NLCrYAaP8GxnQT8iHz
rZHV8F13mj04FhiwO+rsn6Pz0d+FGlZdPEK9rZbKBoNweJzhCxgs+lZTaKs6jKe+hLH1U8AVlypX
Pluyx3bPyruED5pJZy393Y2gwqnCFPeyM3NUdowmQjObnjTXVkY4Gllluauif4VCmWSsHRtCOuO7
IIKgktKmRe5p8wjaEneGT0THhu7yFCAkJblYq03Xb883CxMkFqesRxqjzqWKFvpupmCzll6zxf7j
O1Pd/Xv/QLW6S/NGCvIolIxkVLSvWEt/6Idxn+A1HlJ3F8LSNJhbNBnfB1kaQLaDWH3+9zWiixbF
KSaCwdj+U8O7SlULARVwlMSkBVOTSIHOkrDtwUNi424OlG+dlugMrKePlLHeQ8XaUfompO9vam2z
/uC/mG3qhLB4yxxHkgLZ2AVaFmItu6Me+9ui7pNVPQXQNIzubBFxkHGIixN+PxVv3HG4BghHMpfb
rcFtuXJmO+kYkY/wSPi1QLc6eCM6fc1MwlIaOvZnDfJuLC0P34FsrUnzTu9Z7SiIbqiZ7ILG/dws
MkJqoOvoLt6a5jXqdAFZMNq+EWxxIiS2cIuwHSa1XdEZpDzFVodUZuEqWBpQCIReXmEZLSvCpBQF
ywpe+ILM80vP7Um3JZ690U/NbofzWcbPGfB2tzwwMc9vXc+LBkiFy/NqBqk8g48tWHnvgyvQ030G
gdNOKhWgdpc2meqxIhQP4dJ1S2Lhh40PPiXDudLCJdextXrF4qcDPBwUxyLpryyysiWqAooxEQ23
+GgT6nLeFx4EEq/afN+KIyMTqtiCAJecCP4Gw5KLMYNTp4nl8E8A6GVyEp0j8iR8PSDOCxt0xGBo
Rwwx33t1O4V/Ew7AWRlIWOwsOwKGWQakn8y5W627ZDAjgIymXFSNCUZs4jx1ykD8Ut8FwSd4R5Wn
k+G1/8VhKR67Pxya3SIgVh3n/wp4ea58nkwiMbptoJA3+4rC/kHDA3BQK3p1648HMbC/oGbK0gsl
wX2bmnzr1P/9Z8fCOdEiv63dwVKieArOsIWTYleTu9lA8w1vaSu4rwbEeHUjnF9L1FuCgC6JVXkT
rGKxvSKuJjyJE5sxpIJ45ddP0BJplsRrfzDrcEtdYyZufOMyfOiC5t8b4haclhKX0/ulUy66h+aT
+KaEMYSfWzBemqoUQ6+OsZlRU8dcz3ws5uehiTDwcbhPf3DnIqR1u89KIuFNRj1Q0JS9TXOi88uL
eDZtX++48/8yU65+ghUzrJHfgyybn/tCTcb2PqTKqlfrJ/DgX8Niek4NzkMg/Caz1Kf8ktgu5uXl
Hnit55DtfPOUb4Y++ABChs3b2+Vw2m7L95zAyYUwSGcWjJpwTyeKLjc/c0JglOfRsU76KtxDdJ7o
FJ7qqJmRmIoNrgKJamiBXdlGUxCowba+41qpMcRmmqBbctD2gaDSDR1ZCS7zWdGrGLJw77S/DYJ3
aPBIQ3JA2yC4G/yfnqgrCNRe9CUsa78FC/0In/RVnu1fnV+89gpoTOKSFiFtoQYFFXMeCTSbwyUe
ndp/ConicZQ31kEi+Kov62QehchERbScGGsQIx8BrMui0hNrT6n2QIkTbRU0ItoOhutCVAul/f3n
sQzJY00ZUpUYkRwm8RkLt69tFArEIaz/zpBbe0Jj0LuFSe0xoee7r7koaSqhJp1fHMVitzsgaj5x
po3eWIbzCqZI+bFaVsRRVonHyYgid4hrblPcS3TdQ7chtTzcVPrZ6wUsGNrqhbG+bGCXtdEPWZUK
eGz8rRDFXDvzW8+AYi952gqDwbmB41v7DNgBZmjrxDzjniLfwAS2/mOG5owRc1yLqXOFn5m76yhv
HDky8dZ67b32PiPWQHz56ACBtdn7bGlJARVF5NbnRBGmEmbhMPWYxJSIOQliCHri43wMXMr32KvV
254Ky2z1W0IDG06MG8a/gQpFT/GLpbdMsNkhpll+n3DXW4eN3r1EnZcKYPgJ4wkIz0vB95m4JYY7
rJkusmcZPu96JqUD8k6DYMli/6qUCBWZT+iKi/T5dbX9XAceibNp8YLKyNO0XWHAs1zGi1wZFgKK
6F+XFGm8dRbUgCa4cpYpWQuqr0oSdDXBG9I4b8EfYJdEzRJLpA2RmzMxcldEu5PXDQz/FXIJCmeg
ERd+aYnadmDewe6/kWbe8KLMQGGsPkoZNvUf6xWwWBMKDdnSMPaot2cpPr+mTiV8Wmh7M+cqZJ/L
bQdioas6C8lfielqxfH2VdYRZBJW9NtCgymE2P6tC108BHeVYrOVf7fpeUmEkUBO9sxMjE4c/Cqa
OeDDhahvU4ZOz2CpQ5DrGhXtYdG6Fnr+VZVIQBV9Iox22TJZV4X0JZuAWi9VXzQSxT3ihSoCvQVi
yjEk591/OJLp5h0Lg/PZGsENe1mnrpzllNuDcaZ65OAz0hkuoanMwCPLHbEpcu1oL3SBL+NPzYsB
N7y08SMEH17vmFCS4EEUebE4aPYAQBhklYPiqqP5p6iANQFmd+QpbY/Wq7YOyuGRWBhPXT4+epMW
zx+dFCo/2P24szzP7fNqwGo3OAe30sOaNVK9/3/i2j/wnri+W8lPxv45v538dX0PD8HofDbMCxTR
/+J+CtOPTqbJfd/1z9Fa//qIMIGObWbbqsd99LkrJfPg3GXwPAiXkrztg3GHVLRCP0ZAOS0jFgKm
tXnyVlRY0nbMVZOCgFX/RWhFQCfqAShwkMPKtaiMM8unxMfsSoj0UKVCSJ1zUj9M9eRa6g4dkAQm
V6+IMZq0ZKj71oZIb1rz6tLH781uRROYq471i+4ZoAe9WX2KJoLNBxkFmFJb9MH4vuag4Au2uDIz
UhVgDr8uAfSXmKIMyPBdOLGaQiPOlqogeUsmInOlwnmSS2P9iMhW4QkXgas931jzNWIAS5TmmFHu
MoyXnaSxzXVkHZb5EFIHQMGL1k4dWJ+xE/EnQQuX3c4rTRsR49KV8RhTFhgB85iP/YRWAMCz7NtP
XNqksD6xSwuriGYzn7oZM134x6zpAsCBnMK+mdJzAkiNbZICU6cELGQSPeC9x+Y4RSdEYuQFpRoB
T5SuXuqVx+MKIJRoZtJMNVRaTHBj5KAbkHZwOp5mQiesa2EPXrwYXklH5I+C2zeypcgoyk2bhI9E
9/msYFJKgmS27/9Z2qQ/x7V3deviXada7s98DTCYCUQZ7uWA7xfwrqMe7u39L5q8RbS0vu7m3Nzp
/9gFj90xuHlvfUFho2+IRXOKhBM+rLXZVv+QLGiYThBbYF2zfqPBli68olG0xrUBCgDQL6dSs5yP
/SqfQJxhssVqJqcWW3js2tMw15K1FF615YoxNdYQHyxd5OK8dsxsyCMBSFnbGqpOig6k9g0Piorw
jM5kh4UbiQGDLEZQb8QmP+Vw5GjA+t/6xXugQxluFj6KzloqXNQJWGBeGtye/nvv/W+MSEj/XT3w
F02RBy6CtptC1wOU/RaOls1hmoKnR6BC6VpSdxrqizoBvFF/rzn3Vhvmflg3DfJHjaJIk+BvFhP+
p3iuHSWEUPlIyT8yKGKeqQ+raH48lUEFRMSS7NYRnTe32cEYmpkAAm2U43RWaym1+v6yNZehlCIm
CA2GLPHTuoZuAmWDV3/C6XxFjNr8Y646Iy8d3aE+tVJm/SJ1rWYnqQQ0VyNqnLWv73R50NFRYk1o
bC14HFrNIQd8sgAerviUSx2ysP2QzfyT2vBg+kljVNBXp0QYvMnwTo/UWqDAOU69RmPKUvWwrPH+
U0RKpm522J4Le2rfQA5O2kPe3Woe8bYHU62UAbiRoqB4iZgV8//TFh4vVcK7cx/emokyvR92kBfy
wjEFMSUU5KViKrkvUJA6iaeV6pVnojIiSbrjqa4S9CEYu2tDfY1RfpNzk+3SrqD1ouaPMADFbbfw
mCDtsi5G+Yh4Sj3WWljh2c9duAn/nlymgn5R4uXC5zOZXXD9C8QpcZbywyPWI04CO/GQ6T4yXusN
tTDISCthAoRKLYTlGKNRHsqG7ayTPKGBjOQ0NN66VsIljLQrTVQOuyuRJCBiSItP12hjKZWwmXhv
FgTGqpvMOQSXu+vRZ7OdmDnlJTOTas9ZqTC6ga0FuvnEc90Dr7jg+fkD02w6EebP1czJ24GrZieu
MgipmvdbTjrkdGq6Oham+Zav9fq7LTVudon+GMdvE3WNsUQ9aaiNkXzjBipQsREFktxMezpFjw1I
ul9o9roMtD3ErAHS0Q5bzY8JwfjJfT9tX86G4Y95lWvmycTuEPDy7xC82+48Iuqyok7hoyh9iFSD
5pmrAAkAbqD8AZLFmOaQaaB0BFiXIxBHLPa/ZWVL5P9iA/T9+qmonG0jqE2YWQHEZO5qv6KXxiGd
OCkzgfkgPw5TDrg8XWmfdZukDdQAJT3xhJvS6UNaxUI7C+DSZS8dSuN6PfRZ/5jZ5jhSA0yi9gwT
d8+aT0Fv70H/U0wRrEV0pkUOoYOSCxvTfQ962Q82B5dgyqRNFSfNdl0/EEg32SrASP1UB4W9L6k1
bY26BxMlangr03rnkzMxZP49of7MMiqJF0lCbR0rC10pT3pXXfq3swc+zpMVbMstvF8wrp5TrXwT
88BKXL6m7iMFXSb4QRckS/onkvGquQBDdDjYtzSEhRMN0HhsWukLg8AQ8xGTpOEkqIdZYoS4iFNA
hwQdEKMUmFhn17k+69r94T0gbTWnRl07+EDqVbeUxRKtl4XMY1qB80jAGt/hv5jog/Cerlz6Ybzj
hjbxpJkwIILLcQaRm2knO96+RV3ZSryjXjH2xJVC60hA5Wm5X/oyPGHQUT6/CBUxcZhEUBUiXSx0
LXipWF9wulcXfut+B7QWZDwjWfjvqVlZAJ15E1jIPmCPgpzeNXiRmLk4yaxIlNUqNc/OZUe0CdFq
4UQWXqQB5IQwyEMcAc1prHw/g67ceq5Re6Yo1lqCBeteqT0zrtThR7jQ0N1uuPqCCzPuLGJUv+C2
jkMnKDdaUGPxnVSZ0rQcQfEyOIhuKq6N15Y8Syy+6gX/mjtBUZJcEYTBQs0kx5g8XxkiibwcTwAg
Wl2xHM2riGqClqSu3TnAd6QZt2UGaRdm8+pq0oMrQpytYAGYJAH4Unu09yJ7WR3P4MpDbIUs80Hf
YaeXgPai3SpCKtaUcBLCSrsP4ockFUDIzsgR/On9ik6TJx3nNBuVpeTm4oyxSRO+7XldBk6bZgMP
JlgnTUm4L9YHZ0cLzNnTm2kedVFqaFE1tu4ehG07hQavYuohFZQ8lfMRFAx9541naJOTrmF0Ni9s
9Dfvarv9xYQKdBYcnjshkNqQzxv8ZJzVyyNIsK+xu5IYhyQsciHEHn3d72b43Hh6SHhjhDaCJqGh
xV/2i7FN23pIXLQGDI87gY+pnk/+vyC8prAK61nhYMKPMeJ4qeQFWmSt6RTSRDRnccDgsNErft2R
/KLxE5JCfeEoemoAJubfaTUaMH4MPa5HRoB27kyIPbMFKzvX5IcqrsAL6yBr1qtMadFOqAemlPSA
BrJGjHnmEgVT1dOtk4YNiKG0R6WCDcEMwRDvyiMEe6aEbulU9bYxRwWBaHC3mb5Lh9EIOlEx6yjD
O+fJvnEhS6EkSE79yqP4vFZRQpUP3TR0djeBZ9XBPgdlQQr5j/nT0745VVgFL8aE5eFAOBAlmBwH
8WmHxeuKpbRkHppCGW9wKiKt3I/kWl1krp/oBLC3ibAb2Oxhb/aF1evRqj/brPasB8DUDbNQyTiq
NFZIVbpYK5k6mWx8tkrsHALL9LXQYt3XuGHeVK9JmJvP1ZnxP9bv2El/3k0Ul15YtClFomDMmB+n
M/wPRLX4E5xfGGUJE1jQ9cNgsgOBoFKFsdgCkva53BAZFY2goTksWks+jQUCpT1xMnWymh/D+Pp2
UJhAcgZJIU+b5GKDcIcXNZAqcfGSmw0A3rAMefEBNljGugWQgNQQPEm1h3O6e+JCDy7ONdgQ5x14
pb4UV5N55Iqkus5szH1PnugEf2HZrP34NlIUl6y2tsL/+t3Vc6GnR//XJO9MZ94o9yeh2oL97keP
27aEbBrY7/sxWSLfaJLajYFzMMtTFWX/rWWD9JXZeyIMQKQxeY3TMWfD1xy9V82WLGkff6VRxjFa
oUyj8A/ItZeYNUXk7rRmeAIWe1Qgt0e2NowgHnDOAnDZTso8HZyfFQeeBsUpX3bbkKFVJPJLYi4u
c0u2wuXR6ZqBhFL88Ivlfbjj0TbAKtyEi9Wovvl1w2Ma0APjVADfslfrYSItBIqUzfxzVsN/4W4i
sJ61teNvKpTlPyfh/bXH9jB91d8YTBp68bBZAlglGUss0F+xjuGF2me2pcrMeer+CtCmmru7d2yX
AXCtZNH/3BzkGAForyV/MeuI0IO0qaQ1iai0pzpKX3CM8M2VJpBlIpwp6ZRC5TzodKocmxuorzqZ
MbaV0Fn2zToDKXzXiGPM7FWhb/YkmVL5jkhodupIwAzZLV7dHpk1HP/B8SgeTzNQpfHGMV6TFLQK
W+TSpzYa2/eSlXIg0LePaAf3eKO7/VHGg/O3QQzEKFAWqXJRJfq8cAdnbRc+b2Isi0Q1QGwODd1/
4LN6Cyd7ZkRUibI84rjs+Mryxef/2+5IO0OX+P6SYogEKpgMULcXffMwq04YWMOXNsUG49XUmTv+
sMW8cXxqpIGZCbECFTR2fopPRBK+/FLDZ0dNP0ZJaAwwxlTdEzwqBkuqWVc/GxnoskTJ1kmR/wHI
Md+zIlKeHgR40yIpvznBJekB8/fAXIx1qtYaCKCI88DVg064O+Vap2WM1lVgzbv5aTIrl5wFclGY
texuI2YkLDoMZBlgO7Hwp8/lnhvtZKDmEL6QpOLF0Wiq/lwYJJIoFCMErkR+fx8drwDz8AilBaHg
vzGmls7UPZ1OwbZToE+yQ5xPQrf6nbeyWq15TOwmSzyZuIcElfCCn22k5xUhNhuY2ALXMATgvXQ7
JcMP6YNqJHlWBig2cH8SZr1Oj1Hd/Tf5MdZ7/HlMwGQmLGYFvIsc629BiJI2Hy2WlJnicp87TBNT
/618csVMmdjDSH5nmKT9BE8/i2iavvGdRxkZ4jcQ302gbtOonwQYp1SDEkj8RgMlLQkdgj4wC/i+
kNk0Sv0hZzmSS0JNM/ktqS7MtjN4Gh3lbU/vzAyhTZQZvwfMEZfumAceiCsTlIPQvaGwVNkOPczZ
QpoUTSAgiNfJeY2jETFL7CpMeThVJDRPluZcvIJ9HlZBxbuBlCcnItFobKhSv3iT+hZZ2tW6Ub/6
87O6NGINtbZwypw2smsRgLDepQt0R/tg/JhFWs5KLZVgtxa995YEO4FBdMzEf2lzv2jVowPSPVG3
FWid8M3ISPBgbBFjP+axVs+6opd7CSl44A2hOFNvMsOrddF4E/U6TdcCmwEGWgvBhg7TUE4C1nka
S6RnlwcWoRCSA3Zrtk1TfB03G9iW6+IR/A54ngdimRC6ET/wYlqs8UIVGYxCmjSDtV6CXhABIHPY
LxtCuNkjcHlT0Z0+KhQJd9DeI/8SrdZDv8OaSMWcUbxLDjaLr25AAn65DjfDIebIv2KflblfhRyC
muZUoncppgeBlQqGXqg4uyswjV+dXrDoqrvlUMdg9gCQC4nA7z86nmBfu07QtSmxHKwniCOtgM8o
QfusyWqQJ9ydybEdXRxdWeM71qTveuxnUMf9nAOV8XDYrvHQ6v2ALfgDaU5TKNQObjXoppsVms3r
m6GeJfd53+hWLXjPjnyD6i++ByWYWZbPSczcQ29ac8d2COxEM0OvGX3+pdR8Jv7YU44XkeSWDziE
KA+bj5wd+baFWYsrI9T77RaR/n1yJrf8Wuc2t+hW+LGFpu5KUZh8OkwhG8U/ivMvYpCjfjbE6FPJ
lsvuPQyARFjeiBtJvm6pi5ucMqxJR5rm6T+BVU0NF4HDQpbQ/iFqsgxzxXP0HhOM7FvjR/FigNCq
pEdHgykQ6HrwVRm+3KvkbQP3dU03nidkz2SX4vzE8LNRQzpf+dgWCwViF9BhKUYtrIkNixJjoumW
DILAYhyzpYYrTxDttr7uoBkNEAZlIhyaVvQe5E/NS7fq7mvGUvNMdN8P0BsjOPbvRkYlvc/IuaSk
QBaR1ru28jMuLyjU4ksrHzxSbtPqPKXsO4RB/N39V9qam1Amh+du7xeD0XK6CsW2aZ9GcNxXCMQT
PeqykvZ4Y0/ZB6Ex401jhePS5wsFlBHTFeM4/8H95Ya5gY6wf9AG96rTAmpYojKNx+Ymi0mJTs6g
UQpO5njCHL/7Zm8OxJPaVHZhXk3ilOvR1hWK35AbQz3yUrQknqlZ5jYD1em5mnoFG/weV1E5akSj
KdAJg+st4HiLKSDoVBqqcEd3eY5RB4EsaOkdtu2TuKIebgqcGaV2RIVhl12SIA4bFlfLtWJmK9Yn
/if7DduLwAFKIrs2i9180OjPm5oA3jjCaah4r3f82sxldARz9eGPYQPV7uESkGovQLxFSXq7FatT
nFFeeFfy5WlSmHJGw1zwBcOHRjopLi7Mw3tAC9qwFJYnD6b4hdeuPktGA8VBzzRe4nD5H/82hwoG
QDO3YdgOjjM91RHqf3FmdOG+g1qRdba0Rrb7Q2qOVblU5hz04FX/lLxTFQsNtKVoCe7QKL1Q+VtQ
nSafBkY5xMNzdE9G7pD9CRXjDIG0xDoapufh7up0uzNdXhmDS7UBWd3JEZRuDrFAdc4h1g+jCDtS
jcQkHtUM6OdTu/rKQUsaHVavFWBY7kmmlfaK+FVrgVQ4R//Se8pb/PO6rxJEdmIDtY60Q+GVHhRd
ZdcauQu3jTXlsOJV6ke9BnBZ8D17jFi9tRUnurkx/3SkGUCArT2Tp4VgcioyOtvrtheAvp/sY4wm
PEufInKWY8wUGBp+H8C+tX5USNB2xUTZmq1Fyg7P/K6gYgSLjG/EXHgu8+4U0WgiL9W8Gv6M+7ft
BGbMgFBSRJlb5Gv19X46hUy06OdjaDU/rxN9eVHownJDGOmsFhRcOG+MCMdT8p7wcu1wJyXnbwwI
Cnrrgc4aUNyOn6BAmqVYTrHl33YiPbAwM+fFP8N9RdRZOiT54lu4DJpXObcabgGQBE8imPF2Mz3i
Mq7VQEDH4UIFHU7Gln6UnjGaaMC00oyMfrcVbtUcdgjtsPotslN7bWZo95v+IdikOo57wgiZ5ibB
xy28LQDz9g3wkdrzI5He2zz3prGrYteYN1Mkv/vf2mtqpX6G0uKGS+3CRMz5S6bacnzUC1XiP4U2
x7fn29keALwJQ5cfVtxq+glzsuHmbYClWFw+XbK3gO0bjndTFBsR3+jee4pGJbl6HpJXVSwSztsm
FHw6CfRJadvZv9ddRM03yKgH/kXUO0OlrmCaAAGowQR67MwDT26fYtSubEnGIvSXxsed3OnLZiZL
P84YdvvRiv++HJTxRrNojFfGoNLao/EuxepDJg49Us+HI6zxo89lm1J/GyidXh/rjCFS5XmdwNZx
PVjQkXa/ers6NBugWLsYMj8pUEphy3p6FqgctPhvHXPSr2WxQPBf+DOnvhdf0njJpLTrRU62Zdf1
pItZGBkIAA2pMpsp1PB0TFyf03GFkuEu2fDz43hI8nC+91LqXnquvAD9fCYpEdipkB7qUzs9Jjef
VN71xdTtQPsZMYxOPCw081PizSgjnHthPx+VWDSlbAmISSxGERANxuT/eAwUgkF/HvQftI+3VeWW
XB+P1148kpX4NfiFng9OX+9Ecy7aoz3SaxYUADJkNz1dLrULoYk+e5uON3A1ybRwuqIlk2PypWn/
iBNMOpnh+88/P78PWadF8hKQ3jY3GTptCRGN9GN7IJed28cK/tm0wfG3xMhLDY1C39IsXHY0FycN
zwrPR1GmpATVmmsn0FnQzmqSKGGegRPHZwn3Nz1jS662bRKLnoJ5eAiiLm4HSoghrDPPuL4NRKQc
sD9XTT6iI++1VxQklPZv/aC0ccIKaPL3iq/3Gw76uBXMXaXfdEpiICAAPD3vWsMX5qtbd2q6wfjM
367zYw4e6Ko391tdP6+xWrDfhl0fRvLrHRMxNiqvT2nbwm2dTJ7WbUXYTRAh7HJrDmZL4p8mlKE3
ljY0PwGJW4I0/ww99UhHMbFOTpqLqEloPxuEBzRcnhLC4EaRAElPTlWTRoAF3jUGduEGpnPAkHLt
xqXFAMts1sGwjm6Xr14rHqwJfmvnsKOv3e20NC5Wnju4pFIOB9sTgd8yR3JCl+7Uy/3cFjfflA1g
XXKKGD9K5pI8u+vnNvOd7ye7OLcvmMlH27c7+EpGayXzm8fDRwN05eie/uvIhYeFdQ/umtejgmAm
CQktXYdjF/cbBNBZW/Qd5sOqcRQSTk2KehJ61ilmbYuXn0/X7IqaJWZkCeJjdtsRbL7ZFgfM3SqB
dixRa/D/6acdEpydyr2Vx9AYrir3Gty7Ycd96Il5L/SVSBbYa2HV+3HSp5O8VAT9NyQd5QGud3kZ
/BJMLiRotFLb0hZVZSCta1MsxEcnx1OWD3jSCdexHLT8fdVAw9rDBxCXcrdVBrpxHf/hnA9LHrWV
tfNoSm9LO/F2NrXAXf+V/3EyAXhqu0KhkpBBgWYimJoE20Hag2xmFctfIeU9CPZsH0HmFVHDaa7A
DBwV38ZJ9L+bAJkrCO1eFiqnJ7bF2DHx3n6QZxLNdksUXtZuf7mY2JyL7yQneAi5tZLO0U81F8M3
4QWHvOzcWDkwWld/xvz1WVikOvymwQ7h3b4mw+TB41AYTmgpDGwZeSLR1ji8CIlABZ+62XAfTkqm
ngiP+eOgUSEBik9x91ULNuFWf68hsWO4RtbJr1106LNSWrE7LEvdR7T9vaq2Unqo8KQ9x96l/MDs
xlVzdyC9UkRvPBShztMkFK1MGimX9qIMO4v0ZrmI0D33wiZxBRIl0HgiS0FgZlc6NI3SZ7bX+ziz
gYmFucxarUahE0+1H7Cd6VaGumoXwiSkwxu8MOUhyw0BfW2THPRxUHNHnJF0l9L+7hvsZsgLlfEW
AH5nmWzEOWjLGHvRozSaTUqneKrCbX2bwi+d9Ig9Dis0YI8sJvNt+pY5rHqQ7x4MvVmukeJVNYED
bk6Ywa/JB6lzQj/Rzh+MXqGDMCPXCSDFaP+GHZJls/pNYffyAAa/bGJowzOiU3Nsd4zxRza4s9Mx
2TJi+7zt0uY6zsSsUTg6tsqEOCa8pjhNkg1z5gL5rLhModwdfgPeXGTIW5pX1sxCYKnvlcpU/3f5
UBEytnnjEj96CE0Txt02xJgRZcERDI7ygCqUkzehe2kEUrvHojrGOff5WMZ3lCmUaBDDcnHmkqtS
WYNEBGehT/O9H2EsUdT+mXTVDhMaYkhwRYObVrVa0EPn54Haajh+Z9R4MHNaog/YDHmKtJZVrFmH
L4OndC/U1a5SKFIXgTwr/6V7ouvftx/hRPzKoAKMvIyLiu1q9s9gpqWptIjVzsWLbxoqkiJAtFB5
UWIOmXapcObQS2yPNykblsdOXRgLsocV7ENy2KByxd5aLCv1KUqgiBc2VFhsebPobEdVwLCQ2Opf
UmJUgWdvZJpGp00Kc08mZm/f525Q8+6rLNWgv7amjMqLcYAxPI2hibW9YODKZwYyuqG4LgOoQU/U
cet6m+Z5bFzyFKVLgIsx8cXSv6YwLqQiHCeNIgG7CuXRPxsyefolyHfVzuuab1N5ncQJBpCtA5eB
dSvgMI9v1bry8wNmhVg4aDPLarvuVoL12m6tKr2qxIrtRqi6Vj6Y8aKtYXpbVVZE0P0AITZsS7AF
dZv/zvJLjnhYj8TF3IYpg2gqqvyu0somG9j7wTregmhiTtJb6+8xN4PD6lxx29H3VEUYzl+BgF1s
zRWFlueBgtygjj4XRzqVlHT+J7rF3eJmP4B25RfBXw+R2+A6BP6or2EjFW6fK8W3Q5oIFyUZpRVs
sWjIQEwBv7l+DZ9J1fMYOomV1Pz2fM42xchoPlTNRU0LIeDRgHYDUuqchyxnWANnazDI82L/MlQm
z7Yw3biqzqJG5KagVeDhro58lvW+Ipcv1QH+7Sk7dpAF6cFd5BEikhT8Nflxr4+SQJqbgCgs0A8O
YefmTDrWEaslpweb5CCOXhr49m4zOSt1z6vps7HmZLGExEzCdTrar8pHQ3ve0culfhB0FYWnRx9G
03Jd4S5xHE8FL2hRRpJ5Wjl11W4lETuJQgyjr610qlFwlL3/oGjR6yE1NvZiUykMuvEm0Yb6hNMh
9NRQceWcWTZdlt/Dcvo7EsHsK+dxVRVao/Hbh0ozAB8sFwa2/DNQqDO96Siv9CsuAqH++EhNj1HG
dv7DO1ZiHSM+Vi/R3cIETpUnnP5lOVc+B7ItIivfG0cuacecEf1Xni8sZCTsRoPs8qW5Emsyn9OA
OU9TmaBABJvB8PsQalb6YcMttdiuRSio8yAVhzMSk1pHB3WD3H58h9DoY8NuRUjsGWyYNMmoEYRu
OkK82EcaK32ADzsiF/4TNJt/vTAT+ghduz4KCL3azij5kKcznaQlX5L9Msm0/9NY5BMbSHIKvfv+
oKtmjcoHhmIoLFLFM66nNbY44KNgoNsWyzN+kTHyROg6wQofUxOyK9ZrxBSY+CX/eVXQ5+lVTAyt
8WsNc9SG3Jjgcg3XAzPCn3SNHHW/xVqf/yOlNAGOh0FmZCOZ5AQ84E5VIvptK8cjOBm3M59OPtj8
gKmv4NFZugATBdVp9cgXTkIGk7zfFoxc+BVgdbRduQruFWMeW0ihxlQaho4KM8PL+HsXmLexIVaX
37y4qSyvWmCMr1NkzZXTvdnSg9N7uxdGG0wTHrTxC6kJEpFmvZA1Zj5UMzBRRKboH8oKeupVtgeH
wHu6GKD85fPS0KvWYHKQEtIW6KgSZN9emdGoFwsc70Hi8bLfKjlpjsf4KWj2sHhf025DWdSAQHYk
LRAzofwjjfHT8nfstAf2yTg3FqIXMp7o5mivyAVVJ8X+dK0MBab+jiIRCeC0e6Jn6De0K1T7zc6s
eKIKrnA2DJcYHxgYOS0pVo1Uvm0Tb5JsKOjWq+SULKutxP2OJAzZd0p9FOQxmCgtIMNkKqlF94JP
kAbDjR1EMpvmgHsvPMMEPXhASjvyig+FIa9c6Z0Nya4zxhqeyYGzyIN5E36FWHzjRoNMX6PN9iVF
XCt/EbP2Qj27Tlq6gHIVH+eEEtI3ILLJFfRkJj4/yrmnNGb+zkVPhVsZH7If0KPAHBdXmvUYN2Cp
CnciWNdI8nOGZFQ8xptw7rXKofC8zxpQFhoUnFDHq3P3HWTrQlBUgYw42P0f0K9xEkxEti4Xu1Qy
PtCNjJx69OPGFIdAj0PusVM0FxobZ1ozkAN4yDPS/wsf+W/U0oeBJjrKLyk3OfSrGNOqI5D7txqZ
hNm9P98knXxtLRtRf044eslukdGyim4VaUYqrXdHw1uPzoeyckuH2dw1nD9s/dUrdh/LwewiyYrk
TaDM2dl5qWJLVUkRODiiGYYjoHbsvfBp0bisRxjUoN5zwXNhzLYd7dNDzpUoNBGXqivLE9mYHWIM
7K0WJvDVzNXcWh96zfCkx9Q4fpholswTMEjiaYv4NsFyb3umHUgNAuB4d5q7fmnKMC8+Ae7EipYU
a+QHORhTa94JlKrwwiG1gbDem2VaOH+4efQWPgjVpiw7Wjb61/0LLTNCuF32+4pxbh+A/jJU/uHN
WQNUaKHrQgCrZ3utz5FP39nh1iOic7n5iVcjUmcPHgSyFpeTw8jDa5seH5G7+ghgqsoea2gKFRtM
l7vrTP6Mz5NW6dd8c5RfDySapw6k86y75fUKibJVk9DIFYcq522kfe44mBJLT755JbLbeO5TMXGz
KpEf51Zhy5WewtmzAppAk7rDuMbzl7HzATpZcGY9zk5zQvU9PR8RP7yDQ2ZaBYDd0M8RVyykve7g
G27E+FIODbGP33T4brONgbTcnIn1V9kSUP4DL7J6CY07hLpulZFTaT+G/0Nq24mxcovE4byW9Cr+
NYJPk7d0L2nCff9Wj9oCYHjMH2fw4aA34IsB4sZyVwaVCy8zoy0LxFbx7jcwX/btPqA3XENuqvjY
h9stVnna7lxb8crrrG5h5dToZRyGAkbu/i/aTZ0oPJHfp5FZDbRsgrFBxIFuBD8AyDBA9pUNEWJQ
A+RK325CDlBH5bQfSmP+7rkKzZ++XMX0Zhq9O23xJvue1Q/y25XBi5Bhvo4yrMzHxuulFBGP8rff
yk5qFqOuGVhSQP9asiB1xmjQHQ2N897tuON3FsmLMI8f05qSM2ttHAixIvs0+DKRtN8tTmYcAfB6
sK5F0u/OI+iJzvkZpZlm01wQiGu8FqFx4THENKPbrTvCrcQzqZm6TXqXV6nMnqTMb+lnzAzUDcG1
NrdPBgXfLEuRkXWhSPIWK2XnwNxfoBzQI86b5Up71yv7a51wYOugQipBQKaAEdkQNvBSD57NgcTi
8LQG5f8DVOUOFU9X6jkXKpUitL1lPTd2K7Qg6TLwL4l165iatYXwvIhnOH1e+JuGaVMlnYgZjceO
oPWgLYTBRqPO9Gz+iiGC+djEn8ROQEFzEd07URTtN2ijIMkBZ2zgICqAZSRYVjKyEncQKXlW58rY
udCQ79R+PU8Gm8dPpfYyie7l/3bHHug6+DbT0dwZikbVO0nkAexurCnAoI2elcQm3MqNySpefGUW
Q6xDI6wRn63bT2+pHfuaeMU50EicBTh9stk+LXy+BsEk+fGCnwJp6WKkhFpWJ2A/CC/w4eeJkLy6
lYg6/EXT4lZUasmss1ccozlkusQpA8R8HzFPVvNu8gagWOYa4wdN4S6eV2jaKS19X5+3AVa8f9qo
KtSutX3BMF0GUot1LY68iYxyPDPwpYWpviQZ4nzjKcmToZ9NDl6P1+sg2R5Fto9I+Vte0VXkLHa9
d75B94sz+6jvmMeembGpFLsA8HTAvpnjLVqaztS+KdTyqRt1LGuA8m6nnZAaN+tFaTyoF2/MFSzG
EQlalFZ66uIq0lfsg+su+cZoid1+CLH8mPfOl986J+Nrkuk1pTtBOR9v9Ef4q1ZWHT6u0pWnlady
DytleVF8SWH/RyJEDhyeKsT1cAhl/GIMYhWl1cTvbPd8AtGw5eeEiINOAs1XKrwJ1sAZ5KvzUDCb
GRaHvW8OKlS9KhQPXgcujyPS/0sKzhDo76wgqw8KSSICxLodXD+Q9J/kdSJGJYUvIrP9Wj9VLKXi
XoXzn+EktWw7Zfu9ITRvIyAgQYEKk0+RXysXLf/AOHdfUS0ABOw7QSMaCJu7KkXYwaplESppVSdp
Qjur9FHS0fBYA3V7AHOMLAMcbc2PexwFgicow4tlRlkoD15HhiPRLkJu+xvO5dAQaT7VzEHsLemA
rVfqK3IFg+fR0qBCIFU6dhTX/5KH/Buviq9aiDLI/mvFam3DV2j6fwAc97v9Q8J6mxI5bHiaXn1p
OnTbAr8B519GMaRCnx1VvdcQzKyimfgHm0/X/BCpvvvlHFnwrgyVZY1Gt0PNmnRaVOdprWpvSSby
RURSbjmx48GCuFFYaycAvPdb4G7Ov1MFFlX2TqfDRmSq5Z1A95GoGq/nSi9dOogi4/2dkPeughMy
tft7QKnpr+pSVuBZyWJXJFWlglLf5JBvfuZ+/LDI7e83kSGdIOlVWqOhLnBRXf+T13L4GLnolGoU
Ownc0zRqcZmNTDzs1YkKLvxrHb8LF8XFgFY15wry69GLwW353VTYgk7Wys1H/A5ShM6XGSxp9Xil
r6DRNEc+8Gl7iJIrd4kl/wA2qYKvTA0o8sfziC3krfc7Kr0wKvFXT2JOSwvJCP7mtVyG1WW2uNGm
igw5LFlyVjWozZc2s6Tx04nYpDuLkbfb1+uiKQ2pi9V9xaus27/56Rlnhy99YRRD0x93T3VExLd2
pcwaMXHZ0s/PtjD/LeeQeLsnioHEhsceB5YTpjxtkXFJcED21L9UgGMeWnCf1WSy4g6BPpgJZaSP
4harVbX+r6zKjkNVoSxtgoBpLyGyY93KSVE2ku3hXA0A/Pn0dIb3Uo1S3tLiAwX+gXDnzx3hY4Vt
vAQNdRbOCvVQKYKv3xUOXtSCB/JUYhLfdquCjcIFAR97YSbrUT2I9ZrE+i5uCSOuxVsFP/coGmqV
c5Lxf9G7xZIay5QQP7M4LOuvcJ5ba0hDO2jJvztJxw0UATYHGg20Dboc5eorM3moiSwz7HQXvbnq
azBSfuZlWSCJ+gD8xLN4K8TMV/cBf13jcIsqKbQi3JjQISjMgTj5TEu3w5OTm6qwDmM9VkmmYTpZ
r280I/39J7t39DpHV1xtDLDnj5HzXNPfFRDY1KVkX3CREpyYeKO3KFm6zj1wQiZ0ZR9B6QHng0mk
e0sFNvf8No4qbTrhCobklzvXByUrCPpw4Eeoy1D4GDDLFdURW0DhAyf+fzkWe/9JGwzCucm+3K3n
Ysw4iWxtr2QrrBB/vb+2Lx3iHf+XosDC800fbVqlNNo1GOHICNLXc5wlfn5IDghHW49Uc3Ag1AhW
Cqt68pDKq9lH/rvbS2c84QgJG8MAYqSy+oHYsAkfSCzd+ULYPN5zHCkoN1rNBJdiqcIjmACKJZtz
JjxGZ9T7bZx9mAf70S/cOfdRzXmv1cY6h8CKpkZv9RiOVUyERLoZmKzPTcjeIJcG/iZxsE3EWyD0
hb03z2VwDLEh153m2wMashquxp/fDhPHKjWdEeSg0dQVjCxBdh91xhghiuOHDjSP9y7oNdLV9g9b
i9+jydV6l6a+1j6bEjr3mvRJBPxONUbN+q3QnEXA4D/drIf1XLoWjXW0cosqIcdadNxmIpHk8aE1
bOVJlOKuL4SgCKfC9bshNVV/Uk7Sw+0xvA2lM+oEOj8EL1ISj9m7XWH9u/Ic1o6HUw87jwLXYoO6
QBiZG2W+fsA9Rmkx4QZapbSLsCd2HNh9+MHCKPTqPOm1W8skix0NF6pzqmU/I6nCtQ+7J2eqz0sN
DftaSz8l93aUHgwCW4ap+KcLqAr52p7bL07uGNZCfl7fgPLsVARg5jaJVym9lOpVoq5k9c1K18e0
wvRJuyJA1nLy4SkVYnkz8FmD9i9oMhyxojkR9wxyXI9sdWJeMeZY4NqxrjHdzg/zHfjMPy07jRq7
noptMLgWYDh7vgGj1MpJi0yz2VKgvkJ+DjOlieDr22oL2UdAx3Jv5JMdaya0D27SANgTN6j5ed1I
EAaS7Xhx/HY6pxGwjB5yijnKwwViQfIuSrpp8okrXfNqMK2B2v26KNjLGaQ4GJT8w6lu3qbN2Zng
Vs1e5uCmel2hn2cj2i0nkjRmiDa2+5qYPuUqsQBB5KSW6aTvm7KXkDTR79ofj+iRc+K06oXr1UlR
n8BlMwmiCu1L75hIcEsF9DEN0AW2SyA1DORD8GZqyi/IRnCd3OdGePbb7SLyz6EShj7ucP1t7J00
ZmjF1bNpJUoD1tUd47IucEta5eE69cNnsYsx/KIeeWFJ9it0/fftiXgqcs+gieun0iEl+LOMy4wG
LBEix3m6AUL+1BNcWqlYy6vKSI33nd1bFCaGCToRZn7Q5SuboJnsQeSKiuzlNqmC2jin2tZKuyRh
cAH81dPkY7E/n3vQqCZYGiYiFAFFJ6/Etp0R2r98394Ts5Cls1bch6f6woB0fogu/6mod+UYVMWr
fpuIz7pwNyk+GnUs63YOpiV/q1mhXxJf3f6cfEGZUWBtdIcBfKNVmSh13EJMzaPCWuyHV7x3lJiL
y3/933NeMq40aJo7gpAYrclLG50+pp2QgKl1eLKU927C41HYACuMEhkPS3hudsztfqf+L0Sfd4+Y
mhx2UYbhp/Z9x+8NRFXr/WXS6oZ6EyqH/wcrkQr9eKrCapjbMddF41euhtyek+BUSe0NTzUhbJvA
VCGUdxLp44QoVXe4+9f2CJszJu9RfCao7VPUllnzhjn6c6tHhcr58+SvBJ3ggivHzU1T0Xxi6wlv
786xA9oL3wfhqjgMXWsP7ctG4orvNJrIqjQBS0jPeDPsfSsGlTUuVNYcwPpV8RfDZvm8898tkRo+
2JOEnUrmmyz7GTGRbDHtz5DSlqm8f1ozNTtabCfOyfSx0Ai8aZ+HIP1sPbUYo3vdZd+L6WU0dPH4
akQb0Pp6fvCJ+MWNDpLKCc2ffoB7Af8aMrveKurZ+k4i/+b4P5Ws6/jABwIeZ0eD9WTe8HHVx/PE
e6W8kM3yxpohBN3oeHudNaODMEdsArxPTfHxvzUNC9ZYOVKSLot+1ipQ8EUyG1mtrVs6ZWq3brAI
1NjiFEOSd+xHKs2GmSEdXSHx1kuWvMqk2MbtrQoe+ngHx9lKT0U8Sa8iKnGnsmpzLI7ksXX92XVu
3KB6yUfFBBMIHLUQLNhDjnmxcaMT5oBikyyLTpz1fIjDYsmwPH3OBthc94JEimIccKGdkVHZy1GO
AlWTlUBotqBJWj8s0w09AgV7OXN5KHz7cKhxGWhE5U/O6qVZ5X3JC3bCN67NkBvs+pxbGow+svQ9
Qs2gUzXT3xruYBucsrd1Bup/UYUtvIwCtnSChAOiaJefpasPvyPeJmKCc7rHnoj5iFvGzYVOCY6d
ijAdT2fKTjyTCFQYB5Cx54uNSXXFYvTf1F9V8DT6NBs4oQLLal8ptW1fsiorN+p1OIYEdq1Kjkvv
qiANpXi4JBitNzraHvh+G/msDz+DQHNSNeJ5ihMhf3EZeTCt9R4ZrG96w8t/nX3kIigUCGl4UHeu
sJsYx30Q17XSwwdn6B5e1L+NuD1pS5UIMEuJ5qpOpk03R8VdW9mB71jvUpfRgtAz+8aF4OB6DYyJ
aGpOl5uUd4Sg/NsEOtrYk9vpgoEoWQDlzx7+p4+hq6JPtX7v8GWLAIZ1YhkSeGeeoePTtNDqtP/3
wlLtk5P7JmQUIHmT/VAZJLkauCZAdU+VyOHTMsbZJdV8b5PecTfua0MYTS5C/mL1Ga7aB4pI8b2A
LX7FuVI/9dHPhIqlI6VCpQVVcF6/sumE4Nr6h/LaMARijmds8mZAUgvDR29rB3FMux7KSgzyGKo+
QuXuwb+ueAj5jtPuprEDy+OlXcCpZnwbe7yJijFZfaqWhXDl+CKjQuI2Rja/w6eAH7HyK0WWBp45
/dlMg6QBIqT2Cwkm7z7rUuuR1cvNRz0W8kXyFoIgEKrzLycuJoX3jxAaWN9T1r3+CXVEW4Cvgytw
wNGqdvIzgTkNzToxJDrSMN6BQoCvufPACOXPxCjPaCiiiVa5siWbxMXyQf6v3QwmonyBKAUyisW9
sBG/a2QsG7NoO/1K4kvQrW34O02A5ythzfYCzIieKs3LIXIyTI4ZGyFfKAmsMxfQ3Nmr7ZUjAUC7
RIjgnY2WdbDoSwngKVGVLnBf393DYTVx87qOsqF/XBknmdLhnoUg8G+rQ26w225/kpLfFiiGJVgB
Xm1K7yXfatKA5xURAfea8ZI0rfgRHrjVHKkeHdINFrMCAAlMdnnoWe8QNDdsQACT2LDDDUOs5iJW
E4mMjixZ8eXOjQUkbmALFtbxzf4scKit4WK//o3yMSQu0vYzgNp1QgRkcM82SMQjjPGMTQoK2+aQ
xYL//9hPVCG3YkBLrC3qLNBog89pDSbmkcHQm5EQxpUO+6LjaVIz16FKjD6cy3al6ybdmh+2TvU8
Ac+tloB9O8SUW0UNqKEpe48njmV4sbreh9WQCSX3eX79T5FNKB2YukHxFzt/qwS8Ie0M7xLl5SxR
XghjhVkWboUNvSu94Ptt2SRIM77KKIbevwCi+7gPQL7Ndum/wwnNnVNdKO79reSqlw7sSiDzqk6H
wN4OSdr5lvmjaqs3jgowo+t+2HTXYTti5sDdwGlvyCGtKu1tE5iGwpySswAJmNi5uctuLhLTltrF
Hmm2TPJoC8Ghtx+cBObiRwpIFjTg6sdxgpzVGy6fQzM/iVeU0kfJUCNA9cq/jIqUhSkgMeYXn1Yx
jRPr4EcZbQs0WMjlbOEqRlNLwZnkUVKJWxd6KJKoNyxL4+OBYmLm9rXxx5olGQsVuAlSDl/qaUDU
PCq1FLa/U21UMIrCjqBE1bqoBjnOcf1rR1gTaJTD3gWHvg4MiMnZnLZ1b8/Y/FtchsYuO00RU4Kn
INSbRWKnEdG0wE5W+bgUtyUZQ8hQPCSpN4rWDFKIiYp5NhJdoqybV7igfKtxDdggaEs2vbfKjrKR
AKlv0e8JMU2QZVgQavT0AEs5vS8YrZot41cdYbnImXa/RXacdyboAOvGxRIQ1NB0dNtalibUKvx5
CeDseORhdQVevHMfn8mYcfyxYcgBl8y2bImKK5lYLP85HrqjFM+SFubgWadHrt+vAS7bDWE7D4S6
tYbFvRcJ+BGKDuTaKpmyDaeyHEzxc6eqVan4wdf8fy6ac2EKoHuLUtJSr2QpYPpDBu/vKCjYG+IK
qYuVxUvMg9QoaXUbkTY1KQYuILgMpbmIe7cvUwGnxZH6zDlN77gO1LWcW/KL8orMGrrjaKEkLvol
qjgmGhUoETnWmO96CQuag3pN3OK+lbadWMZOodzfrsPoq+Y6dH9gz9mChwJAKKJYCAid5yU3bAbs
S0FH7vHiScmhMNoL0ru4VmALGj8KtkD801TH/P7/bZmmFhRNnxD0XTwIiOBRPOOrlIl98xzkYbkb
l18ZbQuFezYCAg2AdL2CyFStE9O8lAQXn1SCyy+DLNXE1GoZHFMQaYxqq30FwUIzLI6kjd4LuU/5
B3eSkzUsF8oBYuZrp6ptXu4CwA+8Qr7AwNL0gr0IKVdbEzf5OPDN5Irw5VbbGTY+rPDz6c3+M6L4
GI1X+d/hsXhFRgip7rtdvOon7x0zjOT59f6+9gH7gLvjZV1y34fb/O9wzgF1Ed901NMF32fhaN6F
/iAPcbbj0SYpUKULUy7j2sclRtq9P7oHFJUCpG5j/ON1SbRsO9rKQbz6LP2KwGDcF777qXLA3bfq
9UpUFIhvHYK8mWekkAwjpkttKceibalQOLd4LukVlR62Y013/Nrf78DCWlOw8OiSIlMBLYTPgm9t
nPKwAm2sD+Cf+79mi1RsqQbI5Ygn361OTShtnqXiWnq73mH3wU8jFqxddmTuspSlQPjJhdoIIAS7
Fk1+kCK0XRRuTI7AhFSL5hrWC2I+8GkIaI2o+VfDS7W/EomRZ+wDCicZxUsnw03+DYfL1TmFs1h7
dY6+Yte/vnWM7y0maym3SqXGfdBSF32TYBAdOh4d7BzSHSycue+1XBGp14Ksug6xNxh1Fr1XKx34
jQzG7mT4gzfvmJ9p4MD9oh3Q3ahwoU9lFbJJTRR9fP2v8G4IafJ36Z63jTGqbXITuNeiz6IAKev/
wFE4RQH7xHRJAtvr9DYh+vqBV+/kkvqGp9ctmjfLREE07Bl+0Hbs7NmdQ3JG2hcWt7lfXNkgodd5
+/wCHc/eWkaLvv3MlS5SItQcF2Zk8ThY3wJioJmzBX4HoQJs2pxXGne17DyLuC6mvo0iB1h+j07k
7XeYmxkgn7C+aLdjI4RbIPe2oqtYaDZoDxl3jQpkqqfvV7XCpjyu7WMwuag0eHjg3PqRtFp/KmEM
HwoKZ0lL8b17TLZH8KZT3L8y2K4rHK9cZb2HwwUIa4XOSwt0hddn4GJtR2b5HKIOCisz+9kN/Ckn
0ZGxVWZYi0VNgeydJoK3vd4rkBBKNS7BT+eS8rLC1X7vqCCQefdsCUBd3/Kxv4YON8mHPE31g3Dc
Mwh21OP14Lvf39KEfoMAvk7eSthNhtlMLzaGj1DcjjbxGSr1wx3nb2QKLNGmK1Edic6AaMLOkNND
pElT1dTbCtM83CRMrTRBh+vl0U1/gsXnF4fbFogpt4Sor4vrqUEftL3Vq1B33CWwi5sDtMluwyfM
oFWLbqJUT7u/8RbuCzs7RR/KhWg/5Kt4ec9r1LbseEdZIMmsMGuBcilvYfXzjVCSlsCOF3MDpjQx
AXP+firc1VaJ2nUleTSDsfhdtD/1s+pgu2TNh0RO9nStUMrohVm5rWrSzapjR2NSTa6Q/Ig5LAI/
OJQftoDxAnQgXDhq6OWw5EZl/ykDsrm+jheHNueLEpH1fBAjpumr9fB1xOjzqh5ChOQ2v/cMTpkv
IeIK9Uddaapcx0Cxbzhxtxe+VpBAp+7lFBlFwIFoPKbr3WBO5VlSHLZH5ugNBjNC/ozO+IvSci70
SEGWZw1gzi75chN4GT4GvA1d6evpAYVnuOUqJuWfQfYde3xTKVAIHZQTfOc1M04epzHSbKrVykgT
l881nOF0u+yJ6FgW5JqSBZyz6/LuHz4KgHDKkHrlYZUGjg/q9W9+SDZ2RnXCxG3odyR2wu8QhvS7
WRJJfoi/A0KRiWPLIRQhKV+M/BQIiAaAsWAJlpBhW4X6SPwUO8hZ2MfWWjMtrAMfhZ42FM5VrIYX
IRLg76EVsI6/MiAW3s3SwUVe01+3L6BdjfQ9O11tmbHCEpm7mOb0ibSAFpLQIW7ez9QTq1AckAVF
8zPPjyIWFURzFphr2rKo+gxOz7gocISgTMFEc+3NZA44bLXEz5xt37IZ5Es8OIM+uCCCC8qkM0mi
bhnFjhm4GzopTak17dop33rdpaMfqDHFOFJGaoINTIpK/uvJlvZ/7RqhRHBtifVeRdseBVxn3jJY
DUVAIUgt1cYgnF008ClVsj/Ck6gJw8KEKTE4qPq4V8AI9l9t21izFOYU4MJi3jlOvNGb+fM5x2gz
2WkGLGwA8YeYV8lWCNww38ycH4bQV8d9OwdDdzeI+o6HR0lXSuTdKoY9V79ECOinzRlq2wfubj/P
Kp4vUoZn1Fw6Uk2vrXUncqYmZwJhc3qkfFwLz+ypWvxSXSsUxOeI4DM5+7jcmS9bX5A8D7q+wr5n
MnELoAbtEYD6kUQmuR3RMrAmq0rHlaidh68YlQrY2IRbPFoz2yh16Pl4RMvT9qlm/b4XgTyabBo9
ofrdoPKeY0uj7PHIHcIe3VayqIaTd1wnJBgFw0CtPNyr2ByeBIToIHQb5BVrTfHHhW/KOJc3pt6o
E2XKy+2c6bhEwJyfeg089Bisjtm00Sm4IyNPu85BwB3TgpljrtFIOb9dyRq4UPs/Po6+UTtfE29x
6xGnfRp7PijOFuNT/cXDEhEIxnSikyNkRp/eXuzlVDPNPcp6sX1JlbGdQKSLalvhgzaItFT5FcUt
rZknViVayUmWfWKyJ0IfTklGazlMhjiEPtpzVC+uEr3X2hogPj6/W5lf5RIH5BVdcTC/MBDx7hm/
n4ZJL+3li2ioDsUUKtDEejDq92cHuCOIKOhxdjZaGxy0CWHWowEfPTbk/+Ix2O43x2RAlehYsvxG
gxTwZp+WasdHeRKQFBmRQZAxy/w+OHxng3RCt5NtF8oZ1heIIDZ3Rcnti8NV00bz1e3jLJ0+pGkO
ChIasIY7VEFJvPnI9VnvfrLR0+jaPb6YB03YxOQZj38KQFDFOCeplc3summ1eSWMJ5oWcxbNYs33
Q25W3xqI+V6ssTZZ7fqLgcxv50o0T6gAB579/0pRCprPJVrMY62DmfXXd/bQyw0iTDW3KM9KYFCO
AfFIVsJ9QPx69fuPGz+vDi8XSoNNPo1GU58MXJv/BzqnUVX3soz1incinhCMqnexPZ/otYmR+wzE
Lm7z+AH3o2RqPpilBdJUvJFpmKiqGJbyih/ON3yUkUmuHD7Y/E0qfKCHcXtu++V6K7YWSBI7FPM1
PgnoXXxNSZfEzRloPFHiu5ao+m4MFBrP83n33uA5CbkIP5TQY0N9JVwNsNpAlw11BiSUY/+LjowB
DGsqJYfgbVysg8hc4WxyIpNE73Pe8ZUYXQP2DZ4klF3M4o2zqjky3DkCtu0zFE0vbes8bfN4s6iw
jbOXssPqldO8mVx1Jfe3u24IJ88qDqYEEeePSKvQNtbIXKWO+wK4kEelb3ojZ0CJtniKjj8JOBNI
FtaDG64yLn04JkXtmpR92PjcPSG7Ofqkhb0ZRD63G5T0RjFqfni+ow2lcxErJzJTuwQcBP/AFmAB
Y7LCWLgrHwqDLRcGHTRV72i+G9h3A8J3MTqweuuELjVUBSlcRnaRDayfEjBZcCZxZwxdCyGigspA
B+MtzYHMFoEiT16ltoZ5jL6k1cHNx5aWv5/UVlsDCpPQIcf8H6Cs55Rz5l2k+Z6Y6Tz8EpUP+nmW
HOkcdybcmISd7pr5wuLrOU44334ukqvhKYcgucbQTwfyI6Qr5uKx1bh9z97wS6cvKu42tV5HlTh8
3EyJCOAADHWdWCcc211ktpIHn1MCZUogQGVtLgxK71E5GIPBM5NNZQG9GRBVIF+HOWCbvPA0ARBw
oeJ+aXeBWxyd6KrIbmtH+VGEaZR1bp3Hbq+QRfgbc44J97ZwBhMIIX5OVOXOZv9vPUgzge3YEjMD
4LUlubs4HO28je5ww6k8HMrNOK2qPNCjwMLwaYOLr8iXTS0bb6wTEgowW5Jg8/Zn/+hlIcFv7WWa
u3L/rp3amZsleBjYmngj61cvlObRUhNFotn+ZA3v2/ff0D7YorCguvAXKnY8eKeIoLXxBldO7xE4
cY18Ws9z4kJGmB1wXrgsFYSvKTBR+/VXQo25X9VlXWl6xZg0u4fpf2rc8Ilnw5TQutvAj9UFyOhW
oHpqFtaRd+C0j5gVn3j35j4qwq5Abq+GtxfR1gXv1g2O1C0DYMuM7idAg3/XZLAY1Zb8zBp60fsn
gNgEaaul/g/0a0pw+RexuvKOjHF95tPp0LTi+HCyG4rzU672JChlZ8tSVPN3ndXl0GrUc5Np9KaW
3OmldF0SnC39OJkyCg1pK2sWeoibi/9fOdlD2gaew3mIfKHTKP4JhB8GAEPpf9Qx6dpSFRZ7RM6C
g8bNpO9MrZrg6cpY8k5k1Ycl1aDD8Q1RwLxSEuuiWyneggDOO6QpYv3k2nsLNH8VuvhlstOHlJ25
o3B6NzZsk43B5kQzydZwEVToc5z1z8BX4gnSCL4PK2bP8JcXfLtA6E51rdgQtlrfImzwmMU8w7ZN
cg/4fub5IT07SiHO+0Sj6wsnE0zF5Nel6bSVRqMNxkzulGu5ZmL4YkFESL8PnsdvUkMZi6DOGcgK
4a8YB5J3dqbhmbMjpFFNmauhvRYDZBaZdfNQhrlK2g+SMIQKP8cu+x8Ef3+Ro12tKcDcqmZAzrjT
bmjvnT1bZThTwvPpedSzKxJRoeGrAzaDlE1W9+3i9BjYTA7YAccGpNqRt65Xv8HdwIFLFo5IcGpF
n43DQj3CneMTpYSGhcBdIc/2cXOpVE/cUwuFjJL782Y9ellXvemXT2mJ/iTYeosM00L7hlpYrbwM
ijnrl50ZabuhCQz6sf18FID3GYL5Q3+FHYviNmnF+E2zzeirBBUktljFzYsXVZpI/X3Ds22Wm4pm
E0gEj8E0r+pqVyB8KnM8O5VtH/oMdzzncRGkgC5krc/mwsOoGdaNPqcrGK5eSDgkyJNyDcXo2sVr
C0U+pBHy7oDkgixv0PtHf1ltXon5nXz8C/o9vdscuxre90ji+cfcD+w1FqL/WAqPaWnvZUTuuZd+
vPrtiSJ0cEHwAx2UOOKyRYCSiis/IjVPTQN/6nwAKKr/XDsrIXqGkzNcEGlJ11f9swXLWnypasis
S6znPGrh0R3ePLpLPZVOoRCGdxlBl47lmkl3PK2UX9FV5q99bn+OpdhQ7gB18nBs6xF/0R8JTgyS
9BooKZJ8W/Ap4Pmfe7cCPIe/TjOLG5A/lUghhBltwVu4lkGNqj2cpwxEIkYo5n6ffNG76ST4Yg5v
yQiGi+zTlRFEq8wOSDz+Gl+mn01Xth1CQie0HeU+c+x5RGah75qZKSspQcOqZp8vhLtF25aeLcKO
7yIrbDCagYtcI5HjvNLFKAnTvFPkcapfAstuSpSpEzY1YtQjnWDtdPOZ9MjDeaJb/knURcdRTY1W
yHbFZpTfUcHGLu9xJ5h7yLUqj+R4+r6mL+L5m4Z30J8SkWSzRT/9B/ALdmZ5zyBz5/tGav54rdfY
oW+ZMdL+HIKjyG6EF//0KgT1D1bRaH0akmfBeYd1c2u+zqleyP5aZA2uNg6I9G7jA3Tqlqwk0rtm
YbYAlDXszRu0WZiAAcYy5zfdxAhJ6ODvHjM9hBjYOtadtnMVxqdZKy35jf6gMhnaP41Tc/KxW9W4
RXTIcH3sLyJsRYQLtIkwWU6pihJrWd4eW4bDMyn1BHMaerySBKZnuJOnf3K26xIiT8DcSQxX4pcj
DyZIjyh6GckpBgOb+cv14bkKoOGsPSlvWqjIlLxBQ0Zs01moPW38xh8aqf3JvVQFgDh9+8JchBSq
3zyzUXds4mJSW62H/5Rn/PAfGLoGasojC6cBQeM3Lxl7MMMB1uH+bHwDcuHLr0OJ6gNvlcCPJde8
+fZlVm0yX0trToCdgxNWLW7O1SF58i4hK9f7xdOI28ftKVKScku6GjRc+LgxdyVeNjHKFSj03tlH
CWJ1+/OVdS1qwF6C0WsBg/vN7sRxHZh75xCR0SpUGlZ+djQMpGIqmPkpvYSz0ggtQ3cB5+P/jvZt
sYoUbwpkT6QM9pJZEwjpZRqWdr0eGvvN2lEetdfGdddj+GO4kmxze02JF9azl0laNMu3bGyKs8Ss
9+rqPI307lFHxyObFYF9xqAATnwriaUh0/oUnaisDvfnaKhWRBjCgBxNwuSMCfgSZ8Pz50ShJKxD
kdMK2tN4mBN2EQL6r/lH6JiRbVVtPF8Sa60F0+8C4uSsRcK5xsuODMmYP4oiMnU9Bsxmu5ScvlLS
bP8zfyu0Xo/wQixr6MupvHJM7LJDXhmYvp4buArDrpXfNsMIL4dl/R6FPUTs2djm008caTbK1zNh
1Ig2EE3+pUpqgP0l4WPiRCWWbEUyeZYsOyBC0pyU1uxWiRw1QLUVtHuYa7Qrs5z6bIwdbZ5YfZgK
CwqZ2mDerwUbyxK5+BhHgJjXqPw3mWFosmfGo1G9Y4QZPWSv+csL/RAn8YFF/JdoLszdo5r5Ifzl
b3SrNvz5zXutZ8RQZSEuy8yEm8xFd3fyAjQvydFHkUXzXIAGB5bMWpaH2bjDzikAhpMp82vJpX1L
5QWP01/CPhJfDGPlm2lrncPmoMi9EkPN+w+/nkXKTRNk7Jote7mm5eBQaUZ1mIcxL99HQ2pwECom
/scpkIE519WafCqDUWyWQPqrwCGumzjCO1ZWJAm4OPK9rNwoeMs81PBU4ul5kkv4FlfBrJpDYqjd
55SHdFDcqWxi5KZXhs8UGF1RF5SpsL/vhwbw+3BazWXGVT7wXOkBjA+d26v3Z9z/33U1eB8dtDZW
YjOZUEoxpQZM8tr4yM1UH97j07OuSzLZEPeAj1Gb7ZPEKZKy1OxbpV2vNPjt4klJrHY8HZjhm/5R
uNhgUoeTYWTbqfF9bIUm6GFGuoZFvR3a018NiXDTwy7PASXmtcQ7Hcr4EF/cjK/5y4viOU2SX9OY
ZkR/JGs7G6OQ9O9Ow6Tqgj5PSVGDoCC6Zb9OJJWq9WLyfZrgzJFk+BaHl+rIqiDY/qg8DUPsyfqo
DLNW5gsyTL9/7+oPhLaKiq5jUWTdrbg5XhMCuAYx1CIvoQTBR/5qrUYqIFz/Cyluv7Ll0IDKOocR
oVV/yP8MeB1gW5gOSfoq+JlJ4CTlYNw5/T5DWHhPYVqtTYu46IL863FCb8acirFUXF+6ffgxxxD1
pIYsTfhH4W9IZZvWmHppl2JLcH3hgDcb6Qt206Nu34oGer9M4xB5SkikpSik4ZMQFuV/wYrIhlHk
zZW657gAPZKmptzwTOchtu9KDsSghNA1Osz3+azyDu9oWlT6lbA8X1krIRZddh1AdFln7p1pTkGX
z6GXoD/9HYuo64sFVRunKXNk7BK81oaXTj22iAsd+oP5uo5S4exligo9fr5p8p7EsyilD3j2jHTR
mh8AE5w8txOUjBEKVO7LYLIXFXnFaiksw4fllcLefO/yL1hE7dKnnK/Hi87WPE9jQI+UChN9Wmpj
yu0BVIsr0VxKZJOmSeuyOAJoDT6IGFcoSiBC1lW4w6nU249HSVO0MmWANgyCX6b66iX/knMnfqSv
3PCVqwxhop8uRH9zO05NHCMSlxHef/DfdXo8Q8syHfBAEjtkP2g3t08ZSopFHBCbGSUmw0fVqHkg
Ou8yVwLos0Lb3UYvqYFny5m6n4fjT/7I6f+I9yykwZ9ofGmlinV2MBxFbCjGeRdLHdPGNrXnrz3H
a3B880icggg5rQK88Zc8llXxJfuODGS0k35st40QI+pPIMa/gNL/HOmCaUemkk9O8572Mv4zWS+c
y/lcYDA6m/ze0SeYHxvPREz9RS+WHW03tgArh14MgM3Cg8CWzZoJmVl76m1GOgrk0ppgnVkYDZSX
acEpE3YKA785SXSnmwAqK2jhcMQw4+iY19n4D1l7Oet6l6rYixjZ9wcX7l8UUE5eJHGyiCQWpyt2
+khSe1TodKgOaDg4BSqzmcxrfDzEpVdNGeNW2mUFLu/HGMhoE4t2xPUGhoKrW7nFZzBO7F3WfQnJ
WU4xJM7y1jXXc6EP7PVcXsLzSj8cOXk3PNCugtukPaUs3W3nvO1LHc+A/GSvV3+KClyfAX1CWq0n
Kg+xHq5u/+yxH94DQoydfc/RylMh1adZl/zfl5MY13NZQ6MU72gFXAnodGZIoLsEJmgguLnTYttI
GopYaK+h1vFIVnvXYfYKjCkYz86Htv8UkeB2JhyPHymH+M9qtRk7ZHVRY4Ojn0Jp80Bq/OFSAgbd
CbxVGlhKSqOnrFOrgqIB4x0T54VoGhi5WCfKPJJnKwvNtuIE75fFpoIsU3dIEbIpHFZNka3leE7+
5kVSRacd2Qpdcxqw4C0Zq0bwlHEMirhlTBZtWNIarH02DMuirNAmKZkvGUvEHaO/lNgzQXcBb/94
5YxAeFIvhxEs7Z62KLBxxq8F5uhGdzA14mY0E4zxUy1AkVDWH6wuX7L437GgdDNSI1TLwTpsL3V/
f1nPqUTAYX/b8lGikZF1B9Dxgq4bw45v3h9isIfR/0XmXBeN0+oeP9/wpLerU29fPr8soMD2Suit
s82KnxZQ28B3tNmW6UDaeQFGAM48yfgQjLQcbltm06yQTd2r8M9TCXowb69RI35nigqIhMy8Lgq6
Y41lKzdQRGw/IBcIS3hscse0bj/r1CJiHNqGORyoafqk/CY5ojFwrwAXaxmM7v/21Og79OE8Br1D
iVqhmZRK//n9Fv14YCkcHlR3bHZXlFNutkyGR48BTehWFWdxxdPHPUhymBXUH64BnvpKrD0+ZLNN
cFbUyWLUYpvVEKgrBCfJyMNqg4JWj1wXWt7oRntmYgm3pt5JtN0s2ck+jTGEaL8kVuuocHsJxRKM
e5rhaScdVNsAu4v9lUVHJPBjj1KM2I60PDy4SsPBS1KBMLRMD+InfZkbpH3PJgn5B/t6UfwofeOB
XU+7C8PPpVXSuJ179vWdbC0a49c9B2RayUhTGKd7XJgmd/AdivFvC+d1nJydP3o/uIPCoUduCEj2
vLMEqdoCVmL8jDjtKHUhAkYOby7tTr/qdhhJAxAZ8Gvc4nz/D/XRVlCpmGjULyah/oRIg6I5C94s
6nWhNHmpy2+jwL0I/GBJVjKHIEd5BiZzt0mXknDUns95Iar4RwmGSoZWNVPTueG5vka880Cylf9+
7ugSKv+HETM5ElHnz8TIlTbKSHnho3Nn59/qjyTythNyln2tiQYuf6+TEOeC42vvhwW22C5y0Jub
RVyVoDC4Sc1pC8lTXjpSAKEhF6yHagFlAVg2gLkFEKM/zZteqgG5FOUNbmuIHxk1J6zFoILkffPq
ysORra0xiFXIGiEakuvdsk/2tYXLHwgjuuMwA8xh+sWtK2o80ryDaoEm8OTwe//ki6btnpUYSWhn
ZpktW1E5xY94lpShI5310K2DGehq/zcW8dOZKvR2b/nte0i6VJmWYC+2mOjAIKE1IfxkpWdLDi2k
A++PWPIa6q5QHbQf0S8SZSJb49J/tqivN/kQiRmvz86liGfuG2mkGiPjxO4mCcGXPXsf+Scb10Md
nsgqxDijXvlo/29RbtAxdOEvEMU6vJyFh+jlxQS2ZjNzGitmKGyKzuq5YuxA3xlJ2PVWmMmg1xyD
wkIt/m1juJlkkS5Rctt7pQ1GNCbUHQv72QPHHqwhQsObjdnhKZxUm8n5GgusuWTQVoj2tQfczw+o
9T1VY8mDk3T5MSUjrWLIqd+MZRllkqAZrfm2YwVHcI/YPrMJVov2QhgWu4Ja5ofwg+MpS8cGKFs/
UgsE1HojIbP1F0lwCUYln3xLVmNvc0CfwJb9+CbUN4ESoefdWVjFuBUxM0m5n72Nfl8y/UPIdxUp
d6sAJGlyjPNPDgU0PPJag7j+3Q60x5qCEUAa0jG0NtipV+QjY1XeOOy/EA8cUIbqL7eR4arO7Ljr
FOSh4DlgpW3Gz3bqitrIi3o3eBO1b4y52MXzSu+IRkHiTJ17v5uuXyRl8fRhaJV101Vq9pd9B+/f
a3vFC5UCwVkGWmiJn0AlQSvMvjunAKKj3dlYroyb2RVcU59nPCf8XS0RszRrc2Mvv2eBlRNwH8/8
JDvyd5GNBOnIknMtDeeFYcDe5gvzSzMgOVGMV4zcD7bT+0JiPTORcxyvqDkAckQhxIUsVLVA/VjX
iCigZEDddPwunZbh7YE5XgregrhNkHfuV1FN2NrRJ7Jdg9ERvYU6SyNBJtKR0n5VR6d3gBzCSimh
RcEfEmCPxtDboZx/j5M1JdGeAdPV7U/moNVIJrLcJeu/t3AEacqH9on50jFLY+2YlbdIlkbogAaD
yQFNEVja1N5PHqL7ntbqu0knvhqZlQWSL0NyTOUmxJg1rKd6G/tJkEWTtPLZv2n/Q75UfMoe7PRp
duMKlaQ9sO/B3J2FdnCPPfBq609jeA2PIQAOLYFDKgAu8iA2VK2NDmW7Hnq8qKn5XAKx6UNKZWDD
LP8HNDSnBAu+rvfDkB3ixh4YDijE/vlMBPv5f3fX2oeDy3sRlvzK5REYPOZCc3kLF0ob88vBApKN
EjfE4sEc50scdRwukR5Mx6DOzva5ldPeqrASiHQjLeVzeeDVsZM3BVR1Wkiw1V9gZ+gZyAyGy2Vs
aAewonSQ1A5v7sBDWwhZ/EmG/8HAol3I7YvUA3ePp/L74g1QUpR0qtIbvTRFrZUZF73u1N5QBWNm
d+sWHdiwDsTWJq0U7+R3azfj9fXMghWTUBI+UKOIWWmiDrfeFhLp024gURrqP6iePqECmK2CgClN
CUlr3x41H6orx842FBsUYvRwMp8lA+AnXvSb11tO+zHg1/o0/H3tj/k/LxQ3bwllrg266czSZgo5
BDiLZGVKRf6TKSRP///0hZhwWcENZ5iakBTzyYUJ2onQGfh7rGAzmkFGNlS2fA0X7e5V5CxtucUL
PkSUtyyIdVzN0tR3YK6ORZxARfaYNmt29vuOIgeEHHNBnhSPBwBaZEGpOEMDXKgDiB9gZSVXCmhp
Lkp4QBTSrvn/wXNwcghvmTu5UgGaoFVSO/UJVe4uNeYZSLnBVZ+x7IY1J4pke+8PWss2tpXFYvJc
q8ciUO6YGivRno5KTOL8tplmHbONdiAZWPw5fplIn3jZfUONZKBvUa6Mq8jRjY1q6RrDChGxNQ4Y
0PyuYN4CvmPWZtHZnpD1VruspntosxsmNPm/0ufjrEafAziXgVluMr2mIr5noR085cgwEPWLiZkd
cKHcS9+fDcjqYQqwWuaqW3D3wlzLOFdideBVH2omrMz/0WTf+v0f4TDLN72zR0XbE77sFXnwBx2L
VcJOuGh92DuDMgzzkYd1OOxvGUIcR0wZCxLnfJtic19jiSSR4rpIdsJuw4j0HueE231QyuJLoghE
rWmzhcYp1nIzRFNkggWmrF4YNanxVJDhbY3cXQpacwLkJxspN2RmkWJC8M6NBD4zhkQpzQsDTiVj
Px0b1qKXbJX++ZjlgtfQHhE3q64q8/lJRhs26HTyYGCkiSBcdzLzjO9ow3q9mSlZ5XcGsxx5noOo
t1wFsT7kUSn613kpM9i/310Fd8+B/9h8K61KQA+hXa8pJTNCc6dg61s4EusXOusp0c9pZl5UTc4s
3BX01jMnBg5XFN21wIKOtmANIKCvezJdpwST0sR4mFPMptO2AQJS+/xcCxJv4GMxq0GwKpiU+L3J
2UASip8II2dOGpFCA39ODRiTfZy6a43uAah10sPM1w37U8L2PzRJj2zmrkqivKSbz0YnGyQeeAL8
u6f3WaNEkyB8OyUTzR8z4gSTTwWyzHAdmNCTWsDdb8Ow9jLyOfbxIipnhQL+IVFDLSpTyMBq1KKD
cfPRa5UOd/dkzC/niUUGuLKRzg5BSYFXUrxCpMZkU0S4lPbq97o+3WZQzAQmGzPabuHWifgz0xHP
dyhBPmoTtsdGgbsuynlFCOSLUDF75o97lJ1pDXPLRteW6pRl9GbPDxEAkWuDKWQ/4IbYSnpmLFTf
UhAUJEvLruxoPAmNxH9W0g2sZXL6AblHb+VnNORsvE5ncII4DsqHVtuDjwnSUrHyjlySuMfZYeIs
tSBOffwAAbq4zRkKDsxjUw4jFr6NAbEr8B7b9acqM8MR0XZFO2TdKbHC1CBi4r2tzwkXGbsnY19/
/Xl58rOWEjH/+raqDfhPrrV0e2GnAnPf3NrIQtn/YmWnPyUoZLe3xEll0vyL0uYLDx+X4g+RGqKA
jspbJ6KdZOCGF9egFQStQ0ty73Zl3oi7c0T4BCtJwrc1EgN5e6vVmIm7SXeSfk3fjj3hFjK/rsJ1
JK0fNZkmrvKqQ/UyA8sS07OpHE3WTG2hg0+Mybxm/OHMoqtEhUzsFa7/I8TPoY1nt1LCnsT0tccP
uMpzPd9ojtrxrl4LB4LkVLjCpZgmUSk4G61Dq44tGX3ebBUgJf3H9axSkC48Gu49gG+SpOCbuDoz
CU+tbNKFHpSSJLna14W9RIKpr5wi5Nl77doIwpqs+oRZOnXBiP/s4AhtbDEFhbH7184cNfm+/KVb
KVlKZ8gdC3kxa9npzktBGT8ZddN4koE9z+wRVFD0o7lvnx0mZlGuuR3Eiwar3YMilDR/0jeO65yy
nesa7c/zv6ciAEDE7SnfjZ28OB97afJawzglR3CyFnB9Q9Eujy4JQWVLFzYZhCoeUX9fbeVWk5ui
tzlEPhKMr0q5aRxIoYSVK3HvCzbGwRyyGrCmjDfKUrVLPAtdaAVH+gxjfXh3heQlN0OogdKa6U3B
Rp/4ALL7LQGnfTpdBxWNAMS9FQcXXBBEBk5h5DT9XYt9bUsuoSdCDctZTrSZbsBVefp5NVkH3I89
MooX16ppbysN853f3j1XO1T1V5cZMa/4fxQ5upoWp5Uf8MJUBCytQLF26orRwQx6Z4ms3QIQ4GFJ
H07RJoRYhfFAQF2j2f4Rab7Kn6UbcHiqTmaTyXhUfDLIJxwlgM8F7iT4/z03qEEvZG9wGKdnNkeb
X97yy0srBokE3Ghlt1soMwwawS/IKqAHyl9C96UK9o4nb4ksl4UXVSdnd6j1NzaBItngKKb3BEKb
vV5ruPAWJiuTflSfjkagkYkdG+uRzdC1iuAipI4NYhmgGuUs4l5dwMxw/0OXr+L/aV/W/rIYhYgI
qJykRuOi8lXcY8k9Ya94pHc7KDGVs5n6WK2MZ6M82zFPlJEFqqYn5rAEP7R+Wz17jd2gaOGqolZt
Jzhxqkb7eqg9/vcmWBZtsLbiV2WrNubwXDYWpPLD6dvjV0WwCxbup/LGWHW17jWPeIBmJKd4/sd1
S+E+qsO2FO/Y3YMxUd18AtIujelLfBgeayozFV/N6g3ptRBDVYl+tGu3usIETmK1YSv2XNLB7q2U
hWcl2czaI5ZfIic+SkqAkV7hVl2ABBwC7uNBUrReDXliDDDcs+2atxwS43+cSnAb2jizi0htxtAq
L/VqTSR9t/2WbepMMP6nQmvzCe8XXBBXC75+gMyjO4UOVE2eEZK/vlcLkemGyQdtqgtjCAxvNaWD
bJw3bWdCkBRn8I+hRwgLRydk7O5u8Xci6Xa/HokUEp8Fkwe32vrcMjJSIkykEGyIYboZ9iExbYmv
3nTSne9sP4asVIDKHccK6R8tw31DDpExSQlY0fEFmq/DyLFR0vKXyMPgHN22QC3ZLjNSac/6Z1XF
YMkgkczQktY9DtBcpufAODZ+TPiU670A3nGNei+VWbyVVjt27dmwXN49hSHn0eLf0yUbxOAv1nvr
1i88ezwfkYOTqfqrpk/LYQtgc5AFuRLrfON797USyy56qzRtoS3wJKu3ww+vj+Z0bAxEI3Y07ltz
8mwyO77Lqklj9cY2cqetWHGYEDgj/FTRjwbG3VCLmDy5H9dVFAnxDLT7di9+5fb8rpPIzYCru3Io
YMMD3sX39McoFlg6tGhUr9IKTnafgTSTY1JpTAAGCUfOUe7fADxXVw7kKujjdnwLRDGiYTOnkIuP
Zov6PmVp4ldv2S/QHROsi4XdsPjBEQtNX7wJQhEKcsV1yNWVu6pUqq2lw78s0TBmO77b2GkCM0Bt
fQyX8pbFB0d8F9/74rh1u8cP2YiHXE/WdOdWbzEkcMEJpp8dReirDL7d6X9vIyuBKhsWZmZM3kjs
UeJeAT9JVtAyJ1QqKTncCVm+78p/UCuiptXnIqNzt6/L9OloEVdLsznUX711sr9NEPzdizk9UPd/
ayKITEv8pPZd8+OgwXrMtiajojUsXF6bpEmRq5fxjHSCHwioOCjLduPUbCo1A+CQLfnDXtiJNvg1
e5+jms2FgS2V4T1W0WvueemhfbL4S4hbiif88U91kGmfD6TitE6FnOClpqhgR0Esgdh4LjCVgMtd
sdN80gthk6H9rdET35gb5rpWb+PS4SklPh7/uvpPpFWFEx4RXWADzK+2NRuz4kUrfqea6l+NoBUA
f55cQfA2kQrhL7ZtPBBsRphe5C1ur3SR3kkpfaOcRpJH7lXD8tB8X5uzVO5Vwm6hUsd7/Li1KTrx
7/D9/uLhHuQotfLr42BgXDWsIqkch37wq+JA+hbETpoe3prnpy0gEz2oCHhNJ+ecr6EpERvjYeJk
q9PBaR4J/LSJQprpfvXS1w6j4eLhSEtIIqlGkIdUpLQ8BJjnmSRlVvslZiUYKH48/UpKiRQnXHZB
R5VjeXm1NgENEgPRsrKJkcSuLY1VqMAjF0ANmKJSiMePW64PvraS+rOOWIlL7jOhCpNsNQFa5OeX
/DR+M4oLapnGWPjw6gwjjkXRAeNgyp28pAjcsw2XPyUEbVV7cujJvR6YxZUW2vGwLaCUq3S1fTL+
7x96A8dGkUMUox5LcoHFcb6E8TKc7LykRg0bAFz8dzWQcOgoepokx/xAB09hQQrvBtN/QGVWpbBf
0fH4vEs6GT9WEYTjFaLanX7viLv/JILGg06NvXUrfGYC090yxEM5QARW2crBhNNsz9sSCamCW//T
qP+J1QuDIKh39/Nk6uNtHjTv6pnqZZS58cFKkqCbEzoQy5F1OUYiD9UbLBQvTLBHQTDakUrv6I6j
OspdvNlb1zH9zkS7M4/vkXp4nA3byJhNgRg/xW9SvhYBqCJ44vjjvG95KCUVYPfqqEVezLE0g2ro
ZjJQilAfQz9WjxQVk+Kk3kj0VzIeNP3Og80ZbCpoj7IN5MRdsHOqyzVnenGk3/Epos4bAzeLn6C4
hNXJeNbRJq36vbvtpDqkcgc7VxCay2K3RT0dK8zU7G6zWXMc7b+6PJezwtlXwNZHZCRTCqj2Zmkp
YJ7urEhfAwD0dQ7gN5ILh6bQNBqa5XDvTw/p9WFxKmffzGBxuPgci5nITn4p+tTdgMxNRSx7D4Xs
PhqfOdzye9GZZftGDtluqJVetrhvwoXXL3rdv4a2kWWdoKQr/WVdGy0Vg3hNaL7Bh7oV8b/2WadO
334aqsuwdxOrL03AHdBO5bbApvD1ORM7EqKCJ/x4IwDF7EgzU6G8JT6bH/Klg4LuBjL5JlO8u6Ph
5FNVYfaEMJ6HInxIGzDY2oHE/gFS3l76Gy/v/Oz/LkzIJQe56xMiUQMRpBt/TDX6/3RZSH8v+ZOP
9jygwCkU4v0LsHejMYV2ALqC96Oy7P9T1RU+d3YlH57ZdVBtWWw+AK8FIbhWIbYoHSLobZfxu9Ij
YTw3Az1D7iHgXIVJBFcC+nfkfPMlFvwx9ZfDgtMl/GIe8wusEqn23EsMgaCVVS35CWuuoblLReJM
aHbxNPhAEjSM4cFV6JkjP1SqxAPfJ1UlJOwBhp4FJ4nkpVWaTXdJHqYcbivWNZQlbcHvFOPaxDGL
Cw8MDzGtaE9MLGZLBZaYiixYT6u4no/gh8a0tCg+cp0f7j0iA2rbNeXLz3etFUK9R3efpegONgSO
mDQL16GFVbZvQbhPlNUm6aTVwxXu0aRBXNVzdq1pbVAt+JZ+aZZU2RoxmLSqoyXQZ7MaAS2AkD3U
XIhrsnMee032oePb2phrZhfMT5SoG+kf/wtO7PVS9J2/B5crC2wLaaBmApL7JyqiCNt76a4P4JqR
gKxyXusw4FIsKjLfFWFcf5xKx38aK6od6ztRsxZH5VT0H3VZ7gB+hV6fDxb9NgGhzJzdCr3/QBjC
Ddh38UWDPnggeaXQFL0LtdP9C+ocKffpXypkhG5AC4SAqCusP8uj2nxKo4dmN/MuKsVPe8QYknSx
ryDGgK7Yi8NxvVjxQrPYbVYIjdEMdyA3SiFN1Wp6Ea7ZU+uE2KUuuF8jlAp3+1GcjIOpXDzS0w5m
jQHsd0Hz7i3xjtAFV1xdYw7Q+HHnr3hp4TQPuX2d6uKyyH6SBfeI0k9zgJhyDzitZKZjPkQiY0xs
NAv5kyXyCNqslP4/5t7J8uzd4nt4WtR3KmrOTKXt9ddIfEA3XDuEg0bRaiDVD5uzK2MG1YuyMBBN
nHtwZPgQ+KYBXTNKwLTsFC9zVO1dlyDfLvsWikJpsKocq/g7R3xsWgyCvnveOqul/bwzBIjMhYnP
E/jWogFwr5QfnMzvMtkU+udsAUkc6szadO9RSz+kSEEuf/JfJrx4QG40xsfRRu/Y3iLZAZi/o6xf
LVZ9/cKOMDN2VchhRdHlPo0rAoSmXAncA8Vqo968i7Wbnf0fB6eX9ceB3Oz6h7QaeW/74SqBnYDa
XDLTHjznPSmwhhRlLMktHTGoRFUKkuSqwTTNyEBxZ50IBUyYP3S2MnBYlxvdSRM6RpYufluF2lbF
haBOrfIvqcGQWQQVlm5f6AfE1X3zwiZ9GUNBL3Hgf1Eas0sZA/6syXrXb1smnK1QUvze3UGXdM4K
zJ1vzysTa71mPYk9YJs1OvQAdw15J0pEDSuJR5GJg4jutpX186oJ066PBYXEiQ8+VE5jeJWRHroY
qght3apNuF61b3qmJghpiulTaZF/CM233A9OBE0NQ4zxT5RQl4PzQw1u4jGqaq6amRim6i9YlRcW
edtAg5Cq+8gTY58st4pMIaB5LOmFxVfTPI/IJGWtZERh0UZ4KKuKCyDtOjyHYOLr4JMcC2y85EOO
3DF4izmuwc2VxhXwiE6x6zn7+jwYt/x2Vvlp/COtT/5zg1Ug3gvebzzDqd9qtNRUHyY2NNeyD3Os
lNUugB6vsZGCrNZoojVC9/AYshhTKuQ9jn0ypmsO5u9yBpbeKr+8/4azu+JEnlHLYjHMt93FnD4T
agOqmg4FrUWrtf0WUqgGtMl446B3Q6r/WrYClq+c5yiFzZMJhTWFo0X8ZRC0YB28bSFQVjWeb2WX
U5qr8fbnmOXUewPASs5ciq3Z6594vas4kM5vJilq+WJMhakBvLDR+liGTvj9/mfrKboBKPobCNpr
hr+EO3Jwjn8WDv+rgVhqI5x5d8YmL8lKWFxAvVc2kzO0LXBz3k+5gT3dbt3IbYtZPLXc0SnwK+gz
LCWLHWx90sbx6ahIHCxYxdaEUg1ZdOgMu+6LaYL9aDjcqkGFYmeGbAvpuCKJR85fPX/PEswgkaAF
eXiCzAxoRbo8c9OYT725mWXxyNSw6rrQLxSg1qjGYVMGqKYka/pLzx+pIyk8MvTS5VVyjpZyeRNd
1kRrKb0z/K3rskMiOBv/Uh2StDxxys4kojd+pj9ON26CTHDzbpmEyquLhF41PmM1e9MaC1GAwVis
RiFwJL/r0GsMUBssKB3AEUh7/u203r5mLXwJ6ADXs1ThNh36AQDS/vAfZhwfCs9h8SEAHaeFzsyu
/sT2VGuYEF9N3m1amS7Q9kbnbdSxFxovVDTtj4Msxh89V7rShYl2053ysVNyfgMsPHgCHCU47L7t
W7omB5cHzGhiMJiIbO9cDJdh+vH4/Y9YxYk8MN6ceaeNfVANM6FC0LOY8vM6o0oL0lPKsk8JzydV
tCqxeb1ASEiJUvrPPdA3XbKjGR/9dRmZHUW2IW/cB8kJvWBgrd3VAotf0LqT+Xor/7mc+g0SIeb6
Z5foJaSAocsyn0HVFa8ZmHd2/QSk1QbOA9nqO9WYZXQcTrc2autIFapmvoNGcnbRvsBtartz9vQg
0oOA7phinZKlefss5qfobt8xOhEakbKtPnkWu1Q4f2itKBIN+S8UzpvYTnNl904o/HNluKbXPUCm
dTLNgieM8NAHO5GTcIKPXHdS/rII7emp+KSzwtMFneM+47Re5vvV5dDUqsw4/bVzgT8Buay2q9b7
mTZmdJRvLNE+9q1wcMl0lcAp9TB6zsr4m8QFMR7dVUJvGLGVS7mgXV582Q5zXONsvlK0DJhg6Dba
9a9wIF5Tw+xd42YcMQ2Buu+EcxJyct/FyWXzH1bTCerdPW2n4GeB08Ol+Xu7qlmGx0X/aGrlNIyR
rOg8p6hVKHmG77d4q7Jjhxm5uEVxqyeTwPZHJ4e9Z7Kqvr1Qy6IgseltST5kWBWLhmBxadosoeaT
+WyVvdwFxm48MDLcb7IfK6nGtAVMusQCYRfsC2YqSaZX9ZsW1ivLgOKzgs5gRgPgTej1gvP3SjQy
AsyzWnryQ1X3UVj0Ji6BLufgTOXAp0+JhjXwhonle06DxN5mPYnOUHZ0c4LIL3HiD1DQvb/ZaoBd
U9DRYVXPRrJKZ0igo+bk4Q6av3GYwhAeQhhFpMT4vRD0k7lABga8HTwBJ065PB1vEq2Q+pRlRzEz
udANXbwvjfAzefcHJPLwnasHHjlioEfbt2LX8caGHQjN7zzftHOxEEb5lJxshVsec6N0PRb+TsHA
lVC1xwoiP4nir5eny1eVCYRo8ICTE/loMEsNG8MVlOv912sb984nFcO0/WKiTnD2LLVG4tgWwbY+
CigPCtpaANqbFY2yvIFJHItYCbKuH7sgOAxQM+de7rbMkmSUrQD0jLNexFIqyFyIf6Er10UOOvg8
9q1kX8lZ1TiE7jqq8U7VafV+8gbs7fhtBMXXuoF3dbt0ETXOdwy50Y7DQQCeGcCnyZPO2Tr9yHF+
Z+IpK9peXQOjc7LFh5urUhKgrTxvjE9CcLDHg93d+Jl59ssnoOjqDSsZE+zJCGQqaK4vFW/chmIp
HxNsdHl2+7BrOv+rn5AHZFXgjiTo0BvHvWqwAkatSbacH2t7RrfWSvG8lBaMGaGnkMrDcvnFZxZe
oae6F3gYxE4MzfxxY7gXAMSERqwq0GdYGQIJjKK1TxcguyPY/HdcQ4NOvDuFkVnry14IulFlRlOQ
z3eFa8ZAuNqRoDAnX9cPj8ClOLnMl+2tPPW8a9rzKzpYlj6xUDnxUEYphJv0hVY5gFTGsWkYxMxT
6igvhjhC0+Ma3TMC7A+Gyj4tmzE19QkLLAcFB54v7b73paxzIVNFTC2UuydmmAX6TsZl+UjK+ZNU
T7auJ444GMPaT3b87N5SrCyqeKVQZj5RlvHBtAjd97NAsBd+MFnjl7ZmDiDbsf327PavepCrV24a
pWPOxXoeYd7QW3e5RjYp/wp+vV+IPhRge24RsG6V3VnzfTXwdetCQ6/pYGvsd4mXGunUT06QIn2i
X/z/sqyCTLURBhXD7uFtodKZw5K3Eu8Rl/+lVVFxoVzcWSJWREQf9mQQRBseavlON2JT5j9PNTra
oqQJO0ATTxTAn5r2idGNirGHyIaIpfWEGVCWj+6guYtTcDjiBVNKqCU4+IS+ZXZZJO7twdkAIkxV
PWAJlpleHNMxhYcontS6qgbNLuqnRZuaZk7RMAwnNb9Y9rHVMTXDVylDaHYG3D5RvXS0KVws0igA
Vg1PGw5DgXzRKJ7ax/K/nbfkSuu4Sm7ZOeYYws+7sWV+zpbqzKWzNUV79eaVPprS3rzS7Z9YRkmu
GdtDjAizbusniOSo6yWU7VQbN6PaQ/Q700B55pzPkhxeGqK0mowHMvb3w978tezH2oWGgJRT0Qsb
tPMc3a20INouEHqpvLrz/x4+/ZIrlfkUuvFjHzxDamFmXfrcIAsDWYdaGSZcCIEQClI3wQmsbm38
oUXYTuLLADU+BarG6rFpkOva3GhJJCUoF8hciRkEnZUqKThnZXwb+l7mqPEIV1GG8Qde1kJqDZm/
wLa6XILK1JfqxWswGsInO3ldAJJ11MVnMxbSjnmvpsRG7vOKK4wAqkJbbchOdQ5mdL63vTLyyH3q
5PubWWzejiBhmtc1R7fCucuYoBWSHCmPS98t5hjxdeSNmikXYQ1My4XtY/U1LS7hJSlobECvYj8o
bVgD8LMCpWFDz/Jl3izzNKe6V6/HsBRvCGKdJHyM/M1yCthgRECisvJTGeni4nPePvhuU10uUcQv
+vxRMu/CIUjm78zyWIJF48LETJ9pKepOTb/PfxNoxrAN0dFU+FtCul/CqoDI5Lv8u3YoEfm+/b4l
SKvm4TXAjnJ82eVmxhxsA4lpkmbpJuIFNF4BTEoz6HdnQmW9r33ggKToq3Bi+mgdgT2aTNDs6irc
fJifJID1QG6bxEBmpYLTT4RDxc7dSzjicI5McDud32QgK81Gt+xP0NAPyRhNuIb/ke+l1IbvuGkE
h+PeW76SH4pMEDq48M0O4/JGPVqaJrrGp6DxtP7t7pLQ2xlgDn/MJRWk3IaouF36YkyQGUi2WzGA
CzkTrDtpHVdFkbXO+at3clNNBZbOWzL0zky51tS330g/bBmc3rhoum4X9k7r3RzWK/OvQUamEVsF
Qe0IQZp4D+fHVy1tSOovwqv54GSZmIM2lmy/YL+pm1Ss7nMGbYXCy9Z3N3McEMj9xMDOrYxo5+E6
hM9wFaW8dN+i0j+UbITBrcK7joIB9xM1hiuKtxtIACh0UHyU1gMhPKiy8rqr173EhmE6R64PgmRR
VuAx1UR+9QPYYnt3UwaB2K/+eERl7WGnFlEtnhHEkS3xmm8kHFkqLw+JrGPRlUXgBUGIRFq8tM41
DlTfmP9OqQVHnc0ZmsFNu3/PET3b434ISpYKbWClg5p6JJlH9vH6dN0Rrez+snZpMEbTxfZ7lUgW
jajdCnB8RhrkIs885j6aHwVQQ7px6Tt5jAa1Z4NVbtQaUQuT9SqWWjhYBRw9RYQn1QRmRS8qjHNu
PJsQZmTZ1/O5P1ukqw7pUUdlrJyHt5PMpnxZ/raMtg9z1AJ/vyExZT6XF1k0RNXsJrevqwpHUnwF
VDxZ9S2bHUkiC7FMlGpWalIl5Y8oin5ievynmlo7O5W39rIuZKUxTtwTuVc2TZEvJ7iM1m+YtoH0
pgQksWYJZOkY1BmTtAHihz7JfP1sGBT2GmTEYiFMG2+fAhkz3VJBh5e9BzcoLASpEUjEvBEK+JUv
UEsp7nY9qxE44TbG/842MuaC+ofzl7X/fo/t58t7Vyki3UkEhlGy3UUx5S50kjmJPTav7iPha8c8
u0RSIUhi3l5v0mcJMsuj4QA+WGyCbpL4INO18SnGBxW4rZl3R/BPxlZQ3HMAZ1n/YCdeqwJmQkB1
vbOSTOn3TiS2T8N3YBf0JaaKsE1NNWE6FAmXgZZPDvmGa/DYM7wV3r3oyxmXXRs5lF+Fqb14CSbb
0OhQFQZl2myVkmIPCtfZ3AFxZAL1F09blVeMASo2ZwSVuB70mwq1A98otYMJ9GyRyTc5Nn/IZrw3
g80vTB4/+yy9YdFb7UNSUwgM6QodQnp7P1tCwwy23g9hOQX+PZb3UmrgYtUd1rtp6MgmjZJBgyxl
GuilwXrauEVBCrBPG4rpzHXXEuEbIFv013P0u+2FTFji0o8z1GSbzIfJ5jZXqv1x5HjOwa3GQuAl
xb2G7UvG3465dcFG4v+ltWXJAGxy66K4HZvQyFffY8r7rHGe4GXZl1XG7jK77L4klmhGhUpBsugr
TjbSoqkNLICP67d4ftLxp+eyZt4MCp/dhKw76ZStnngA0mZDAzYmhdOnKpT0NbGJzKP6M+PpB6k0
Oy2BavXJ7l8Fttf6f79uUwFOjY07QLgotntiUL09Kdf1EBKE3Bqs2cDcR8rSQLg+KYF0PgMDPVF9
jE8iv9tyhZp1JgMFV9yCtDoP0mhcHnwYzDcV1a4RyX3Gx/o0rhSpsKn9rg4d74aXQ0yA6ptTw0od
G4+cEWoPNrllVLis5l8XB87OI7l+XIvmI9HZfpBO+x4n+G4YOpKJvip0xr29Q5A48sOme0+YhEME
Bmv+h7nhJrZhsUVkaVgjWUdgmt9bJZGIQY593gpOw267tjP+XhaDydE43RkGS6lkJ0rnZMyy1F7w
s1IWEYa0VyRJEMpZtREc0YQeWQKOSio4fOqtREfekSyIRhnuz6AJ9uemAmntTAsihVleHjUKfoYU
aSG2KBMwTzOaFCHkxBuuPyURJhtxqZGq0efm7TrSGru36+K0KtRP0TTPTmHOeVWohgoxE6ZW88b7
QGjlQMuwSYcQmvD7MP6wTk9xhqA6QBSk6Pd1/Almk2P/SQRNROwmH87Cvp1y357GEc88aCGawTmd
MufPjE9Awnl6jigTBgXBbUtqWbhn0xX3UbHBMdUGO9AV9dxiVbsOnebDYFmbc8VGpXTDgCzNXT/q
D0DySuCvmq9VbAdTbKKF+m9VlFIMdRXx/Ev5xWQCTTfhIijWLaEovxRE8RwNuV8ytSLeE5J6ZQcW
tzx8Wb9qukyioVplwFg+Y+yEXQTyYiOZx54KA8xF9xBM1A8jQgqaNFh7YnWgvuCKij4MHp/G9USl
cagFOgBzgj3YtZx5pS6zYdmlTNgAR7/HA5nQblhrgD51TC6KDDMs1cd4G3GODNNjMgQ2iBQ6LNQB
sbnLx8YZDmvr53ip4MW+A0oCjgaz53au6PlINRQwlOT+dvlIr2moomBgKdmcO36BYfR5Xv67HsyU
xC1uvGwurPTRmdWtWRrHMc9NErr6bDJyJWlOSZ3pwHDrnv+P3sskqquusJx6/lQYa+5z9ouJeJY5
UWSsvMIR6FIahder1vkhGlUogAjunmaBc1f2tSZgdkN8WltfM5hkb0t1ZwrRMmGgkOJCD+wgO1ij
V9Dg+yeLLxQf74+HHQGSdIjAJ1RI6X/KD4JH676r06o2ganmA4WoAarxPGBEO7jfvKoi5fHsM43H
zu6usvR2kFHkOchHJP2lTZi4j3p/rbDzCta6LjxRAimY7RTkPR36EDisy+Pe8QM5a0CQ1d2DFa06
CGI0BCJESBRwSP+y8yQmeIxGnZZ8gb2optoZVdkRJJOP4Z+z9tVFicenzm8L85XzR4RYVvopTFsL
+p2Pxgqzn56WOq+y7ck1/AlqYpEDdI7f6cn15/jpYgmA2JOyg0CF8xJEm7fysxmv+DKgeewk9ML/
WPwsMRahoFsni4WkvIN4UAC3Be509ebxSCGM79t19cty4lF9euWBf/kZIP3Eux8XRb+Rg1utRF8Y
4cZ+jqarnkyWbNM4lyLWJUtJU69nuXUYAtcCaerLYt4AOshzXS5SlVu2ewJIxotEsAJ3CRiNt96h
PlrIBXSC9L9JRSYwxX7CZnRR1uE28bipiUyZGVUwR7k69tTQgfA5mt2l7chPtu2AuqbEh8KzqSsP
QWnlHOG65Nk5eCE9BGxznfAL8QetQYU0K4cnlcME0UxRnUKncJo+yNYWu9J5FQMZq9CU+xSt4dj2
su/oxISEwdoqhv+XJZKKM/Ep1ahRZc9I37GVzxl3gAwhoK0CFi87MmYxqv4auV+X4TAVXGvB6cwP
pYt2SgcCf0aoIdTgdY032FEbLIR65Em88/ROJDud9l22GW9Ryo9+VqhpWWRPudmr3LPXT4vMDLiE
MZRTLICsLXeyDZbjapD9hoo3FTB/fBfaKjfBY2QPuBg9zsDqT50bxuG2G+DF/A6RKpJ5DbMY6TL8
CVbskTBWAkMgpS2uDxC0e82otjbqwANFS9/6c8dD/Fe48QYFxxvKQTdFHQPePyw17LQR/fyZxsxZ
26POOSeko22cVopWPIkLfSD9d6GMSHWDD5i4pTT2hZYY28TAiFeKTZy5IqkeTsOFeZIM91u6VSkx
hfOWpNHGRNfRAKKApYlandmRql9acf8Yhj6Me119RenJqoMksN3nHg4+hK8QWUBJl935Bi03/em+
aQk9rWDlypsL+TQjI3oYQXGeM2N24WY1zEpvl48Oq4H8XRyocadVlDDfThKe5Hp0W8ZZv6mgD2hj
55c9N7OxNKpK5+Ukwo3RVBP8Gh1NpcZamNt01J9M5a3HGEzjVO3KwCJKXpuNqsZUnI5C7PNv451Z
6LS5PvZ7bo5lSMZiXVdMrvY1WAASMPpd07k6Ry+w9bD3Eta+yqMFiujeTDzzIfRdK0SormuASzmK
wtem6cw4q5uZSiJljXXJmaLfvLhPP+H/xzRTxeIuvRzV7u+bST3UDKeTMm6GjfzadLTWGimWhZfz
eu4tBM2i7RmfWYtmOaWZh/QHlgMHf2APpt8QZXTxiv0fovYHCZcOPiNrE3u42u5BHjUWqJ58Eucl
F4XEdFyCNRgJgu6FSTCifq1c6Skx40aRzSJhYP7g4Mj893mFiDOzKqiDz4v5a1hcD2X2JFcfUjwr
+kbMOU7gyicC3DUbxNHAZAHICsYCTVsqI/PuBQE8EYFutj9/aUaJOx0XiWNxcsiwMR57YsRvdCsh
SKAZGmvt8q9hKopvyrn/yREVjYDzRe/Chx8ZEKaMZGXQcpqHB5GlGmTEAsiQk0YB8YNNlmq8VjBk
bdqrUCc+fb6M5CFax6Fq3cK5X2giS9IRqG4rjR0Clb1fbZQCe7eDUUGRkGeNN6wzbzmRhL3w+FYg
Kax4jYXujeVZBBQvKd1/w5PWsYUPHm1961G4pIXQapIRDELY79VtD8oVC3CYfc+UBxc2O6N8Q+JO
cCfN1tIdTZq2HXzUqTMXfndSIuHLbZn8Q/94QG/b/59B0sFEzxdZ9JJN7x8m7vWL8xl9Ycu+A0Mj
Uex0NyZMw7KavxAEfa2qae6Fl3ir70rwpTcHspEz6AG0w4sza0KlZBe9XEBmxWhoyNoKH/JyQ5cK
NUKAIE3X0G+vMOFermsK43NZmWwSxY02MoIkukWDkpAcoRxJ7ONWp2zgSH3qEBLFV4i8Td/Chekz
yagNESb+Fk2j9f5V3AWHY4E0FG9GjloByCJyJNGwxDB1mVS+j7//WgONPnNXKxh3WXXYO8V9VEge
Qlt7G5UHJsSVWuOj6+edBS8z/phqp+KGaITjChDps5llswOsZ+3BqThJBV1eaUmE7YN1RrjOn5ik
bHuTJzWfVcZ3RAoW+7r/N6QniD8YH9sPO4T3cpjSbCylO0H+lAkpxXxe+oQFAke5oNweMRafs8pm
5d2ii/UBm9hSfL35hGJCQbBLx3jxt0IHhr+O75fMUyMi2eO/C7dwBXK17X6+LT4OjkfaOjLboIKv
vU+H1fj1HHNK+HHXpBezgmfHtA3nwodKZBB6UsPlkbuXmTNHilDpohzvjpv4wyGLbin4ecyZPWWq
32wjfGIUHNtmqMXWqKoEr3bzzUXHZaQwo6kGMf5iz7vBKq2TFjTduQeqjxSRnLHsEKqE8OTGQI8Q
sN7lNBGhw4o7taAzF+VVB5Qm2Z8uAnbLOvt83VnkM3xZ69iRyOyoXVFrV+t3k2osRZHyAWeKzasQ
t+p9FQSVenJosFYu2pLSIC0+/33JZYlqVX6t+tQUFydN7frkANdpJq6Y8ptEh9l41yv7qIy7EgtA
ZEVTOolCCTOwkAm9moVXZnngPZFq71+1tvrr+7KTVCQIOZq719Fr9dWrMe4lZjqq6eiJ7rLH/5vy
lXuHjWaPcAhA9jMGCh/xsj82SKWJQ0nbwV/Gk60Jbj4Ta5+TArWFmpgYI7xhdAobsxa2dEgxx3HS
5vuI+kkimCN9VZPuqsSrfAoUzfN4BP2vbY8U9YGHbsyEqy9UcFwUeYFVDXXEaYzBJQg4E+6Ebcp2
/c0/YmXUjr00xAT9jO+r4PDShQaxSbp9FwKHzKNVSIHrXNVfoZW/ozMoAMt4sVm+51Zxi6jWSkr6
x8G4Yn4JsboF8vHsLpV/U8XKWwDvFzbyIWhFGizrO5Q9iOaFMvyWaabaec6sl/bVhQjPiK0XunFj
1vVjWCyWnv+yJPV2nmxTaD8rWJuqqdiYsrZpKPKG2NsJylbEDAhkBjt5zsingxgCoy9R+b3k+D3g
nCgBRwd0KJ1gX8ABFXNmpPJsAD5cyg4hg5zdGFiqm3YwtsrYZcmrOvdZjulHOf3HRwRgEv522+Xs
ZMSCxDzqxc38Lpvp0KwOeG0X2QtRcIdszzH1ZkFzbGPGQmPatad5uGIpAh24xzDADdazZM7EMyt0
xTmCBOqd1XoTqZOsZgNJWAVWJye7bE8q7DgIorcCqMDSSwBdmyVuz00ToXCV8toVYEE0qyn3CEIx
ChKB2UREU9PfEdhZyNxI6xsgYsJ5N92ApWgpzgfEvnFYBLV6dLOxfItykRqLakPPvM0Vr2lBb3Fn
kroWWVgcrhFQiUSxrAuW67LuE5g64f/2GVvGwndxRhSLauj/4sceQAyRYh/ceEBBb1DlT3wO1uFB
BcvKpAnXsQEsK50189urAlZw9Ve0YdiPA5bf0MeaXSso4R/X3R1VTdRnOx7qqrx5vTlMo7rWpDKA
pD0bzQkGJTwaBSB//mMj4ElDtqJVL+Tszo971isLMd6wQy+qfnYzdZF8c5gVFpe2ULc/ZlGazQS5
Z5fg7iXz4r4boGTpgX5pDZsMhO1ZFYhQRd+nFbPwn1YwYcvptLfm4bxmC6EOKPDAnq7JkrW1635x
sw5Vwy/PtayumoH7eUhCXbP0E3Ew9v0/OS5x+01WKDMVBMyiXDjZ6vjQtrRVBAsrDCdVfhRjaPP9
HP/rbJ+38Y4fIqiMbRlqRgAoawd1Ht+DVyNrYoESlgNi+VyCGPmMzO365ja+SQfDvRYrqT00YBaU
be3VfIU+WQD7qhSvuLHeWv+pXbhCtyuRZraTIzSvns5X0QX4qyqcBGPdiOFqszlrZog/3pww37Az
q4XpWDNQzQRc+YPHMRK3UZ7DwGtjS/42k8mZeZH2hbFhG6y49FKcuI/F6wxfRCqJd2Q6LddLnjaO
/6V4OjOja1Pxl9ogjKHxK8eWg0j4wmtdiijmpVIQ3ekSvqHk8aSa92IwVNgSKcoIyVC98MhBeRJJ
bEdawpD5BXiBaNuXmD0qG8I+4mXboz81vvOgROxy52C0hhIGTLXJ9AbSCY8IdkbBzMiEUEC5sv1S
zqEVXiwaGMeIwEBxFUrTKpA+17gvN8WHHYW0erml97E6ROfyJOOLwwsg3zFoq0R1BDkEvUiMrFvI
9UoqAHLl4Nz9jQHiJ4ofiP1tw5oxG/kiEJz61UTBJpOa12AgTcQaK5gQDGGE/8EaH7SAR0QR2CQX
dmXMToKYzx4wiNS9E7ktMs5Ea+lpZsqc4N+MqTUMfWu+vouRKu8XDy+gwKKn+ykqog+N4Og2Erdu
88xxrVlIFKoS2po1aEcnHpoDQDdKW0490NYFPUTRLbi7NQJjaD3A7baPTgyJFQMX9xpv7l2/+kbK
R5efYvvaA4HTTckKal1d0PfVPGiIPaOl+xLJ0fhHK7gz154d0F/iyyIl+vaof5cu6hWd20QoXYWw
bsJZVPQbXG+ofHvn8TRQGdWwFbE8+7wj0zJCfj6tpSWTwNBPWMM5kf2H3CX1j6e+gUJltrhEMAje
E62pCXCnrTxweqb6DU7BEeaCkBfnjVw29WgjVFen9TM3g1VThr58GeXTrhacdfZ5fyVbKZcfonB4
5FEQO9G4d6lv/EHx6nI5Yr//CAXVk4bVuHQjQIDNv4e2iW/9Ax0V5V6aAi63J2ptUHhkPNxS0LNX
+HouNI4BVJUQW8fzXnEyWJwmwYgIMXDU3PoCRKLSBBZvBRyoaT5eJbZ/BmqWIVl8972Zl9ZJBgri
N/WiXvhmYqCAE2qG/m22KwjM/roMI7YVy6YGDBumic4vhkdJMj/eEATBPU6l7NzuFyZYI7QS9jls
fSgL/wbJhLVz9FNUzjcwPn1FYyMsa/NUYV4/Zpb4j9R5JPdX0g/Ph5+ZIt+ql5tCaNrsxc2i3yw9
2M5NKRrLYR/ju1Tb6Wn/wM3SioLKwWD0vse2ASLK9dr9SEkqXL7V5KCNkZ1JdQd7Pgbua9IGZ5EJ
uazyUyoWxmiSJN0+o4vtskYUcuEF3WViGDaujkonThmSVaLg4wLR2SBb0H4zIyFJh5z8XKc2QItx
1Pq0Ey8ej6rvBnHIcsNFg/T8EruyEBHzB9bqTk0LxR9HzxjgbpPjHptNbMZowUX7FJsQvoRokvcH
EPiCQHe4AGl2u5sU4Dw9fWj6vIJcR0PCbLiEX/XXcMaW6aeWzX7qREG8WMpTQZhi9epsHkYbzLP6
ENVKetbp9+XzEGLPRDsJZqj1rayMqpdcNWYMVolVG2gwpPRACoFefhm5k9s+t35UhQzSE4zoWVOz
YOZmTeurR8zD57xdYmkNIddW3Eu4mnMH7YtHvr/pn66EPmvFTojOz2eS7C+p+82AK8X+9sVsvHRV
11pgUfvZ2MscvqKo0zAd4a3u9N+GwdXtut/whN3dVpVJziuwGPsWYdxqlvrGHWXsB/T7AeiZlDxp
U394X1yliWoSDRLE8ruZxgbBUObd5GQfs4GX5ivPMLnPQbIdERtbglBxrnLSj+oczWY6YUDsRP2l
y4M+RLIKvGouwBaLucZaoLlg3d60tSkHwtktV7uhFS1jWXTQ6wwOZmoBoYb4SJaWKLmAVpd/h3u5
WnPU5oeN5esKxyRmGUyVTs+Zi33HgUEKuJYpKM5qhGPW6u4v0J98XN9G5VpZPt06b98egeWzYcY8
rXZPGKp1kisvXFLhKxXCHgRQO7exxw1A3TZY80a5aCWA12MJCiY/G8k6ww6GHp2NzNWpDqp/Qyfu
2H/XG9E7R5N9/cATYl2jpK+9crYQttOY2I4J/3/GT9n4PUFdc1/bKiTrN3PBMGQ7iP6gUMDoIq0t
qawWr+vKewMNHYsnJs2axQsRT0lVUNlIm7tdSMGYwF+sXGmYx0XStDO3psxNeXpxyFLTue2cKhdS
6jf19tWAuYxMbWsAgtrDaL/Y8PD5UkMIH/5Ei9R6uOjiXVbU+0JYdBb1yQ5wX2Lunt5AkrjR6KBW
mNm9juyBnE1cIwEU/HUjLYfeLqzHuBpADVMyknnoSqWC4rONOXvdziIqU/z5ISXBEfvXy/0bzBaR
A2horKk3RvBUqF41+zbMnwJ3GLPDB2R3lZ3EjxI4daz9l5gtAe0m50YlPABHiORBjxUrIo0EBCoY
Z1spF/uRQDD+VBn3UZgfJIBrbbVD6GTvAx8xX1sEWU/WGlKI5sadSBVNqFXv94/Pkp24+cavHYZd
YkExw2pJIyEQNI7eDPEZZF67MOYGz6iGg0EGHt6ejZrFsgLquPQ0ACRXAX1qw8n72ijxKEVNjr7D
n8XS5KSHoJ3FOKxVd6Ww20lrlcZUjbu+7hS5OuU9t4P1CT0AlAp90kQDmUiy/4FLtXfn75xbcEij
x7xtZGBH0Q9S4+c1qmHXBNmlgCD+nB2ikPjQd7TefcJuabxv3nkwBdeWEQ+AlwtuFGoCbxqdtp7w
I34xipzVAyECDkE0nxxqb4zq8uZjfuvRIwbHtP8pwCITIbTMytHoC1G+0Wy+dNEmvWQ5j1mCfSK4
D7/x8F2JXLztOHKobZNEBUA+yx7/iQb04LKzB/f5H4cR1+Ez41Z1hKz7vR23qyK37+mHSeZu7Uee
6HeNen3pnpsRkm5qUK2lPt+khgb4Rw1cvbJ+GfuG2favIBtx+myy6o7z/1p4+oJ3IWqicb8J4CWy
7k1YoPBAoR2KZFzJSYrocRWRq+P/NQDMRh6VZ1NtwMHqCzqLvLkLSUPD8tbjDnM5L+pdLq0XQZfw
0XJO2ZXM7h2XPHSDTt1zw8+PUW4Gt8uilZXdD52lWW8Mpd0NcuppTUBPuvGk4CP1FSP1PzFjjsvu
G+UrElccRJj6LAUV0WuF1tYif1ATWSxzhIptrumY/rO4LiEaNBbZ5Q7CG29Lz4n2Xhhk87Re89Pj
2YAQMeY3Mc/HdDh4D9iceXnr567WZrerj7K4QlYwxh3DX+jXvsVEllXw60fzk3Ohop//6eZEJFLd
ffX2o083e6xoHwdKlUP9VblK//uP4yVzuJWDOVXCC1mM9c5OWoa17UFOZx+wMu8prOo5eWhvj6D+
4SLDAFO3q8oeSBFQ7YgJ117n0L/Lc7Wyml2DRhw8MJ9fyzGIZRB90Uzzsp1bCbfWOjx/RybXwNi2
KEklNtPi+MlvO6wGYGLRxSn5xzT9MtGQm4eEhtNITpl7cSn1nakSS92ph72oDNJzBt6tXz9ERQEj
yKAV5K/ofXXBB0pJbEnHSGmCBEZHDh/2ESpWOUsO+gtNzcGO5+/jLlOqMjUZLHTfSkqY6epbwM/i
nOwZGyPEB+OQnqnOnmRomLohdyUBhZsUV85y9vLOCuKgKMNGiapXHBKC41wtJaHfUZKMamf6AIa4
1pfGV2JbIrSK4sIHSSUjfLiT3ms5GsRL4x4s44IQthyAtCtpPoq0MD+mKuV/gSZhnNgD9EeWRX8V
nJbTzeqnVp75qlC/LvMZcp+M/WWT4GCdkOGK8/S8CaN0xw+/9K84ndlZ/St1D9jzmMpF8Y7/HwyH
WBvFuSHdYsV86/Cpc+mIRalOik+TzsbdfqLP0APVdUfJhwfAJrH6KY0+pTWS8en9Na0M/F0Cg2j/
MaNkTbH16fcLGY+/64BLrcHJnfWQ3811ixtr3vokd12+D8mCj4acW/sGGRQCigPBgL085TIBHqhl
nbZ9BmcsgOMVeylo5zpqCtHP7E4xcuCMxzsWizfPqatHjeSysmOAhEUus4e9f5JFRc6vIi9vYItx
RRd2kOm2EI/LtWNeOU3+vC06QuDN2qmW3tFeD+SKfWU71311tEqNDzgKO9y685eKCLOBKreTP3NE
RWJtXw/gG0JJTbTyaTqxgEfA3pql1J1ztAUOFoxoOCtyL+Seow2shRChqMTnRjc594Iklvy9h3QO
20/nL9CIB+y8qR/NivwZEGA1UtspO81L9VRpepFq5HuoXk2G6JB+66VTqEfkxfw90qsNdneDUolZ
j8q/7akO/0G2PGtd9ciy5Yd1W7SRRVodyXr99vXfLtgFeDky/cmebTvdb9RIPLur4fHIY2lK5Wrn
qpMywyBQwuT6Pb3hLU2yZib9Ggs7PcBJVzZYUy8SYlwXb8NsYjTdcd/4r774C35KtHHaSC3eiAI0
ScoiIBiNf6O8Pa+ZDs9Pcl1WdGLRMO8bfpUSaTAEYa9bLs/EGDCSUuX64psk3eDBzBRNnITChnfV
G5DLPlQy8EAwXFqw5qyCsQ8L4RFSVKkmkbIRAOBTluNfNep2B0eiSprYT0vW+BKfXQuS2Ou/HwBE
fu45twkT164YEKaGRmOijOehNv/kDY1V+l7DROpdBFxoxYSeNclbrtSSjf+fO11FWeGx84jInB+r
jVF8/ccJvMKb1S52zESZT1f/XETR/aY0ln3ecn1AG23tPPwJIMIDoDNdQ3vU54oBC29OtjWBdZfX
dvCYtjDX34YC9ElCx49e0M1R+M6LvcdtwTqi2QcLCBGCf+blPk/pBpw4NZa/4QBsJ1CLJQpP7XGu
o2kDWBEZFnt5Gj+TyJjg9pJrkN0hdiJRoQ6aP+iU5WNr6D2qa/0+5YjVL4vxSkgxnQYYF6uEhvzd
hpeL2pCFbt554RyhPvFTb/IOrZmaiq2zkLmqMss/bhHRFH9UcRsP4LoAoDU3ciKyYTzhcRU70AnF
FLICzfWqPNrQus0YIlASaFZAIbhsLJy0UWmwgMlC7iTT+/ESAdR7O1E+R2M/MnXMWNpwzC81xW+a
Zf4PGwz6PuGfvBei4A+TXsA8I4uCxYUbnknXngTwOf7qNSlEyzMn9ar5DkFZL/as0qH/eYG26jML
Dhp2fHi4F6XRm+IVEAWUa3wYNEKB+GNEWLh6XJwjmVsT7fjjGkLmvCup8xDYnzHT7OSDh85Ari6Z
R3SgAWyTnUTdrGEnv2/BbgqNwxl7Oz3RMKJLnsU2Oll1i/loxYfcr6IzgTGxp6QlmRUBoZhF/D6t
mIONK7xXdFrtXZqPMQe0pMY4N4UE5ZNFYmMTOA0F3DCVC4fF2HaCiLQCJAP7N40JsEZh3e9EAQ61
yHeWj3NY+bOLPudS31c6FFFOpaTyVBhTUc6gCeOMtIka2FctKN0YdJLSNEZ13Uoue5cNJZHYW1Re
4/mqWBHb4I5MuQffibE4Nj5ncruQk2l4sZCHp8aYM4T24N3G9MmhDzp4To6xll1pXBv+ygrgr7gt
C190b3arPTMvnH5t5MizmqpoAyZ3vvlIGvGJioEChxFTp536G+hbK7xTGmLneTTSL63BKtJ1GINV
pZuLqRr7C+pFhL+ooCqp2hJWMRxKwAWKdYcRA/xIYEiVg9qJXBfSLiaP+Psv19iECkr/+1iASFWo
O7a2YcBWhCfcyphRwZy/YiA6NQXWwbnPFY63I4KMp7XJhpmcJ7dwWj8A3oxJMAoxEYjAHNb8en9j
10f4sIMEg5tKgp9dQu5L+K1uSpfw6gjJ9OQo4ssDBvorJluiZyjDhcKSdarlmIrYKN80kQ5P9uUO
a/n16a351w+wYJtJ+H9ZPfMFMx4JhQnFkivPAvPMBjUK2S7o6ngw9qOosLHS5Soe3LUF2Dmi3VWX
drE/x8lO5mHXn2/3C17N7Wu2B89IzbdKD4BgJoEQzHZGP/QxOEsZf5fNzLNyPHagvkUu6P/u0/RG
OWoyItNNY992xLlbgRSlSriacLY4TsOq1bgYBLPTuF/DDKDBD28xFeDFCLpYvvnqoWILjDWuxO31
3X5VMMaz1yLBN9TqIIU/eFra/Z/rhvNW5Uht7FDlujsCfcj4eUMOoJfEgzrqDUwn1WUVrCLiCF8x
ay+aATQuGx26MnobkbJQn/NourN6tRwGkf8W01djc3WxC00CgnqF46NXcd1APvPi2NvoHejRW6u8
u81VkrRW7XKi06kJJQz07k08Zclj7OB8qxrUw1B11ldBQTFBduuXdHGwrXz/QPhyOSua3Inucn4H
PzB2+5JyizKh0FZYcnqrCXTzIquVpb416A7cnz0fwmv1tQlL/bJytNdl3dJwYPmd20POf23qcmUF
Y4+vMCl1Apy9TWsw0Fdwv0QCiwZoREuV5Y5IEhIJYt7pTQlOE3PrNpN1QJvCOwt9uGBCWMTS/dTs
ZAa2YvD98PA3xijfa4gQ50U16jSECz+9ok1OW0rrno2rfaDLg9V0IE9raDxElS4AecbYFG7HnQ3I
7nRl2J5YqEKtmVzYNkUhrXOfcRq3qMdbqG8S2Gbt0CKQEn0OlkwKHv+FV1T7eUhNfP3L4DY8jleJ
okhA3mDdHhHmXGRW5DweV0ToP4B6latCZ4RJlqj81eWk/wMc+0cIpvjGdbrUVafyOuXfusQfflxE
ytaLuV1ICSHDl8qs9ijguwSTQOlhxZjU44Uje2B0ljYDSTJNSI/BqFoszD5wFEFDmoYtxSiI3Ajq
gyV03F115A/D2cxg7XqbrV/NycBcLd2pj/fFmmkqJF2xxvXjzq+8+2CWJPUPCA8JKPU0+O1lwtMK
kgu6CD/vcpVDzyLgedGYaN3wD9oZJfTIohY9Pd8XLoCjv75RK+k4he+om0aqHGh55Unx4UnudHGZ
3beSUCowC8MLklsqq8zHeTOSbrO+d2iF/XDDz1v6xX5eLmFFKMmai7L90f9RYngvkLK6wXlLkPSw
16bzE652B134lIWvEHsUM70gf7KByyYQYzCT7TkWvoRAl8KK7+cMqj2Bkhsm/IcjGH7c9fFtr4Yf
2N7v3JLNb/aONTvqVZ1wm9A0yhr/4Lw92wPGfGB2xR5c199Ls013PrAFkEoVUWJ2Dmz9ZabuNnfP
jmYAFXc8cbGdJ/M+yv/01vA6B4a7H1qfPZfXw0cs95qiEzl7vpljCmqB92QWHYbMNfRp9nvgIn+t
P7HBo/5RuG0gmSlYpJsF2AFfbO3ZOSOB0MKq+fh+R08mSh3632kuM/ZeePVNuNLhSlKbAySBrP7K
9fgFE5FTO6ZE2qBOoL1zKjWiQE+3s5kvllwsAuXa4wXF/PtParYqThDaSCsWC3uu1uwr8SGgHit9
H5VX0Fo3yZrfCVVNgKXYLSUfGY4krqQUB2kdG8qHpw4XvYwTZtFpzJI6VRoZFIc5bybDhaqP7VhZ
oaLbuC9clek5LFV5KLXCv7GeDSCL8rNDSSSqggNkn/9Rf9htnB4Q2FBVJJJOkNquIH1E7zteksN7
xsQmAZCYq/eRCgJYxz+YTEEccjkHLNm8ymo3hyHoKQG+EkXXB0vzEXVwaJWcDwofW1VuxFrVHjHV
0Ec9O3a9cS75wNd2J6gGTBj5nTywp2VvHcAGGEZANRD0+aXXe16eaTQ4gKYA5E4d7/2/KXw+lsBX
fbDW7SDMQi28DA79LUy5Uo+qg4RkXYT6f1+W5ygR2VHO7lLHwgc8Fij5oBC4n+D78gXwi707ssWB
L5n6pgcC/f1wVfyea6mpNlGI3cqRU+TOTsGB4KBMpeSwxen2nbJzhcalxN4t6/3h8+CbPpLbiGlO
pybIYHnbkoyHB8df5gRjHIqQP1FsKsXnL0YxFYp1GXTsh5CDdAq5ZCQyy3iBUDOqA5c8GRdUOXKn
ircVRnFULCs3OwHi40ff+hO2pH1CpWfCFD/zG8/EfC3ldfzwa/81cotwXSufxShTVc+yLm9pcb+n
Zb2M8oMO7oOPfAP5RX/Cld6naEwTb11DINSXqTXekAsGIDeu+JdLpPKAk7kch9Ltf+udgSVHNOvW
HeD1ZHw1p9/8WMJP8HgVxrYRYrWh8z0VSwZ8f7BZXl8EJj6/ffssGlSxQvvMzjbzZoeJSV98s7+9
/DXX76iDM1c9G6SS/m+tVXoKPYFF2YppQHNlgddoqoOJCxwQwbz3vOL+Xu1hxsHHQuwlsNJfsHv7
xsZ7T7f7dRoYGW68o1iMTrw1Y3RfT+A0HMeyamY4oSYVHXXdqND2sy/RRjpRWN8WhXXHJOkjYxOD
6coh6xFi2YM5p8JRywTTWLfrTpwHW2iCzoXxC6fKxtqdxtaE3Ll0yW4XOihpTE7J0nEkVEbumA43
Xq6fAUs43QZODWN7heAwBRGaH01Hk9FZi9RAyqk4nCei3FAKVoSPPxsA6NRNy3z+Y5Q+Tb/B7UIr
FjfnCJwWQPresMeTnt6tMlsRmaZJVyd4Yv153TIkkGflYSSlEb+Eugp2Ik/xzTQtpugpMsYqWG8k
yC7ZDaDVQvDORuEHR3VlNSx7Yk9go3sWInmRbXvSP33qSjDJ5gycIeMhROrKQwBvdsW+nLE25xw/
e6LghgUcRQipcPJYWH81rmHFTMnANCsTdBVfLFVqAW8TcbmeU13g6xeB4//j3bV4v6jGFvP2EcBR
8lvlVo0BX3ImdHeFscae74rDkW8ED+wX7l54mEaWBG5uylhI4+zR16QoHUwKKaAHTrhyoymDVIo6
0+dEl5kUONi7O3HyA4AHcpwdHc3xM+OFlZm+bgd5htbUnRIlYAyC/0++OtP6UJD61yP29nr8l7+w
e9rcEM1aJsg9rZ3TitOVU7z2ev8aV2oSDvYtZZPK/Fk9oLjNz9TQRynoS3fLgmcCug0uW2/7bLcy
aOFg9eCrCDrLCf/W6J7FqyKAnVr0yrXd0+3ZtVrvuk4D4JuMvX5ua8YJBDOZEkt8lGKIdkkr/0z6
nOXD3NUq1b071G+03j/vyaIeDkxJa/NQ7/i1RgjcTvloeDh2ZuEHnUlAW6yWNcqxhl25JaYTSHrr
QlRMKpvNcYdg9i2xuG2JrMDFOMK7VQGqxJnd060vVWNKQfcb0xlJGJTbuYy5xAQEJyEYNVluFvFS
UhLnI0I7RCtkIF32T5m8KLWrlxsNhDYL72lABh37z0BvBnM01YoAcTaOSpNzEgiO4YziEzHSPih7
wY2FSyt334ZxrXWQ5GBJArIdM+vXdlmXZVcc/Yxho+v+TnWpvPJOoa3Nj0+bt4cs5lpEcXPP2hvi
/fDHUnT6ZNUjkAEnY0Mc2rhofDe06+NSM86UfqfMxO4x4oqgcS571aXbCGB9BsAWaK1xMD62iMeb
vxqEXsrmtPz2RIzVv2WQzwMZsg9dFMiI0ZhkdeDIc/+OKl8ZiSNItZnTMeU1mHv8CN5d8nTNF5qf
Fny9ka1dlhQU36qVCXpk3zh50zaU86rI+An5ilksjznR+jm8Wafimcf9kbUcRAUMyPZaqIG1SIX0
tbROJV5SV+iWWFXkMAOLDJOXbDVYc6P1k1SvGLRA0CTBccm462LpyBeFwsRDFnT74xZLuK2+BBRL
pUC4bC+LlGlLJ/VW/S0vbFdgeG0/uS7AEP8YefxoEaJCL5DaJrzWk0A8R6xvoWSN9/cLlHMpyreZ
EuQpDpEkz5aWBIt32IESorzbzLoH3GKB67ptKqRcFyFQCqIGLeurtDUspq7He/6TlNYqtY4FDVgh
BGbRf0/9f53h6+sHppp4lG96l0CfSqa82B708N4xdnTBGsApdJhnC8hFIp9HiXp9cQ3GYTfpFJOI
YyfWNNkEPbk+CBIZCM0rcnU++mOHaJ5YwGXUiwLhK+hZAp9z2kVp8A2AZNKD5+4/pS1kB2ku74Yt
E+as95aMBu0tZIIhpoQ+IQrVX902Gpe05wOWpGzsOUkqAPIZ2s+5yDKNkJbczpvSgws4jyvA7zUK
BHmiGU9UgK9OzUiQjEfat/FHPwpW0FbIPb8SYUh+HMpJ4nE/8wuF/8c8lJx4XOYJECsOFyCMrv/J
Hwwu0IjD8+CJM2hTTB3bUjBT7Vmb02Xm8M7n0ijekKpqtxaH5LqttbLonFOz7qkxUCCjAHPXb9XC
JgW1DPENqwouUQNcZ6MKOu7o1Ja4PZGYoF4od+5uqfutyB2hrhjDspvPhMO6R2JW6wYhQAZep/ug
URoImVuLfVo1N5p0LuJsurajZvMTUY/wNMrJHLauxJPSYS9BcSOGIojFEonFXEJru66IfY7AVdca
5Q671VTA3lI94BhMTwjovxS9AJGBBYIo9Gn6ZunBpRNIvvPWg6czushkxTZ+tk0hq6Ct3ow8AH1Y
+Q0rnkDS3mPdCVT4dYw6YqYvReGsUMY+gpZb9zCykX10s/dX8dDWo+KGMn3NHTLUylq/jAyTiM6J
OktzeR9kOYxtkw9I5HPGJ4/xBIC2ob9e4toweWEOnjZDDBrfjLyph6VrGZkBbQXX77N6FhYPyDL1
LlNPdpuhsDNkbPN94zCvI9B1ea4gLeCF6QbSWq3cn11zWw3vZ3DAYXcMOtuTRjo1BQX1GhoVf8ux
geLS+RdiWzq6BN0NAbtdlR7PRpGVe8GDPHHkqVlsUVcySVV+2F82pNkVTPLLarMKmebieYclJMzq
Sxas7P7w6+WYJHIDwy6oObDazUegMPK0il/NnxcFduZyP8FpUfRNJDKDtq/WbDwwWAi/NMahPqyd
gsVY7MPDmew4zsD9yR3Z5NtwjPj0yphFHXBo7yrPbZ4weRgz+VrF4h5driUmbRjRPOdGQUbxOZFn
MuJ0naCChhSUOyu3VxdBSw9X5CQLBv3/m+cy3BSVyIcp1p5vuvEN1Pw/S3lA3TpIupFDUG8dojue
/D02axK0hU0BbFoTY4nSyRqM93UxH54mBFRfTbaYMKuytinRZwq7z/5pFV6iY9OegSfDz1YUMhMY
6JI8tWIBGcRhJYAteTqyiSaBR1enJzqXWlEppeM6XUvTeZ+uXa0rRhp8LbFg5Uu8B16e/LED/Nrd
Fh0z4SAU0CfQFNv/rwNdicd1kl+SdNgT8PkwB0CS3ng1FhN7bGxmM87yCVOgYUWiHTkGKMJ5OcqQ
BFtdozuhxLnMTPX66qr2Wa2/i8ZxmWkNXhSCJei8qAKB2yozD7IH/XtcvBCzn81Tv/PDqMOTuRlK
OZdXCxHNkD54xwHG2yQ77k8rHsCL42lfd43nBp7afKrMu9EBE3HDNVNiwHnjbUz2GmFjZ/qj5ae5
HdYf2MV28knguH/wcTVB8+9fI0ZVyAUP++LoALfZDi9ykDwB2dP95Nj1pfql1zU2i5vxwANskHn3
PMly8RIodLpS5CEYAzJj+QPcwJ6cmXxgK6S5dc52pjvYQv9mUtCGeWuKsjSzmHrCb7Etm4tZHdH8
VE3uJi7SOq36Mc9Yz6/6rlyE/tN3kSlfp6FTgPTKekkcTHoyyYlOcK+4+uoK6aUbA3TTppNd88pH
hAv0TtmzOGuao+GJKsH206J0Mxe03yAhTmA8OXPl66EKw2ZVGl7G/VEy6MjRdZsUh0uo5MQFOIKB
g8mPSLMeq9EE+BkITUv3LzmzMnfcgT9f9HB+8mn+Qk5wSdYs8twR2zHXh18b8a8f3hg05PsX+Haw
/BaoPLifAwA7FUTlNVbCacSJB2kf57KqWCUlcyN9bTZbq+0ljtHRFsajCXOEU6sE9d84CPgimtDH
Rfiq4YfPxvAsLFk+ULX1Yg+XhyV9VbqQQlG69g7XIGauNk1Jibe2hqTleBREEC6qXF/pG/9FZpXF
OYLsuXeo4ECmf1auvPs3BGEaggqrljJ1d8JwCcCYpEZuzB3M5MXz84z/tCD0vOSPSIZNmG3Hy6Kn
nejcEZXzjKkL+tCQNOQkb0X4Eyvm9ZgxZhLJz+dGYMEb9ut8DxaUOcIvCwA2uBiO98p2Eb7zOdWa
jVSmDf5sVQwXo0uR46/b+zKmjIM5mrMc1audz6yHy0eUPlKlagKIxUO0WdpiJ9GbAT/wq0P4Odt6
dJzCNRMMexDby2otjuoAzsq8nXTPMJpshpz59rAATLydpnncvl8ESafmh9pf6M70dV3QLgdSEuJi
bchCBVa+bUvEzd41kiNWDFv5JCwNAMidvl2MwRdXTzJe4n0my/ghzM8sOWfTXc1ZQOw7q+pZBYqa
/RzNlu2VAjj/LbFrt24bEA63A9eIX41z7QWcxzoC5rPBQ4gpE3lqtZppW54h/8eHV3GAfO8P1leI
NUJ9FqEuMTw+a314YpjcVkvrTQIZKk2XIST+mlh88dGk5iifltB4QuzUHjUqO5zt8GyIjeTpPOKu
5+W60iriMJn2UVxDXMBNy1fdgxIevmlSLr0T9sc/8MaNm5v9ofYmr1TbqgGTZJtGiKtQ5TIZI/Rw
2JePg3hFpNuWCn1UFGa4M1GBt1ZqhT6ZgygBC6HIJPILo3Jz8W4lMVY6J4fqJBntlj/wG1D+wJT6
WxEWdTCS7WJV5BvT7teaydlm7kqqLX1K0tu+I0a8A1Vrw9k4A480SR1u5Tk/dLr5peS0TYChModt
QUyqIO/SafycPMakmdIvwKEFETapYqrF8VlbXGX0Fr3rlrnbyV6VmxNdpyGgoWTIQfIkvPfW26o6
gtHvae2Xj84o75sQf7t8OLNqYt9qEaZgKO8EJE+Qs60aUBr3Uid4w5sVUtXqyRFiQPGXgwfnJgXb
1sCIeuTbd3kYTmQZ9Vaz0Jnu1A9WYk8z1JNye6KAFrs2JOYVxEsuMex7EEnTB5cALSFm4pMWvPwf
SF5narYhL4KkgeSGFpCYcI/Y9fX8GNSUUB5AaE+hRPuX3ruwMwG7ydc5eOLCw7ozkEAAtYZYs+92
Zc722/zP5Wd//A3EJhqcO2uErRsCxzbfKYr2bfR9Uf34pURVfuIjP2rou/os19aGNOJe2phK7095
Z/OyRM/SXRAHeiStC5BU1v9OH8UDP4IMhynf/LAOYVDljDEgK60yIoFdG1dFB1n7Qq12mp+8c6Uc
DjrBasFQJA/b2imGNog2plOIZHCHghcWr7NRvc6YP9hJaCi4GETV+WRUmAgLe4SBdeXnhKF4TCKQ
eGOC4PthRgMlOQbWp/C8TX7QKDtugibWWHip9pqg1pHVM+vVN4f+CfJb+jrbIvi27cbMi3pOOj/H
2q4R77e/gHI0dcs9bY/r0J3bEcy+X1N7feQMNozzKbrfdFWNyV2b/KKa4ial+uIhsc3Ni407ivnR
B+BRZyh45d0nG2F/lZOPH70UICgvECR/HPhyaO6slujAX+/EoVwy2o9dWB0dCQZvLkWrGb1bSkS9
8TAP+F/GHBhZGjrwCCk4Tw/5I/tRK1AIbC2hsjxiPizO7fOv+fyzZjgVqtilSs4cPPFl/CU1sGhh
+43cDgYtGfx3QJWOQV0y8x4vbC43f4qDIjLWyOno9b1NpKw7lgRn2+J8lcVSewT3HKPrfBBZBBgM
FP2f3ss59yS6qZEKn8eses7zLRNALfCNqxRNp5g2gfVCoBeNvz1A97/xHkkfnbxUm3j3SW5u46++
LFPkWJjpVDjvDAqHlx/BrE9QdZqdpG8HFwgxhZZ9l0v8RBN6JPrSAm+jcgEeqsrYGcIT1sMo4fzF
/+p5hX4Y9HoRYsZ8XAe0o2XmKCcpyW1hf9BhIT9wP6gAoFZyqBExuKg1D+nFFmkXiCROHgemo2zp
xt98RN+nI1Yj97U+q0U5eUT3vJ/WhWE2NtRXBtZHofh7qPz2G6PZAPD0Lu/2ws14x7ll4BrzdcCN
28Q/fR3f6LnvCrOVmi3OG1Bhr8RW1m3DFQsyWtPOf+7tozsoYKocVFoO8UuJLBKmdzTQ2AMZLjaV
TL+zJVxHUoHiraceaA7O3HtgrJM8M0zXNx0TWfv2PpD39L6MS6c9K+cYcaYaRpGdOWtLbifhaeK9
vSGOITLM1N1p4bFSlhiba4+9y9g8JYtpARwd8e8fXFYAMfYGKDelcjQAkEA/qVIRkum8LGMmJ8Bv
790pislX4bG8B6X9rzzxmlM19HSClI+f+QCpp+MQ6L7gYzZM9ER9BZ3l6W/lH6Mj16zY8IZ6+/hQ
pNFL5EsumEBwyiIxwSG+ME4mDO43EGD0n9fNhGUBgtBjjBo91YlxQp+M2POS+Y129vjLZXQ4EA20
TCdqKH8yRRon4YT/fOH1kPIZbeWxy0nHUswPOYn1M8YQPrrDU8IdpxBgZf47xz/emwp6/XQq5Ge3
WBZkvQi/oJU/uMgSCGjurCXn28GIhTq9Akuhj0FWIzImpx+NYjh+aFUIcKDc56lV2G10shcwftri
3fYvNR3AqAXpP8x3/zW9C/MGQ4LGK5Yc+PnZFom5oFko92iZXGjfUm7rtmMQIdhmrd/ZEZEsI2QX
ErZ9LSYAdvqMll9TCm1MM4hudl3PK0uL3IbS6gt8jnzJp2uyvrxQLRz9uHpMBvElnCu+dNPHOU04
UK9V9KIT1mqWjvWb/ebgvv7RDOUkRIGNOWB9sW4lo0XWTJzykaRqYYquGQcLJlejyKPSqgxzYsWo
we/RXZ1HNPUb1lZRJS9Q0l79EVqA4sb5wqHU+sItLM+ICgkmXh1jeRDP7vZpzn7msnDvhxtvXyOz
GWhfj5LTVGr3XswQ0nFJzNFfR6p8E8W96cu75FzNj8xIbP71ODVfxwFW9DDzbBuqbH23+sA0e/Li
WYhnqQh1alOCEbksTmUHpJdlUuwzEmpMY+eFYgeyVI0G663jJb5VxPrC/SkBqvORyeOy6qCH2F1Z
EISD/JqZAGZ5o4C5NvKs/Bj1vsWQ6Zf3gkAmrfkiGxj8T4p0ouFu2G177z0pIXsWvZtGautFsedi
kn6fgBlxoDUEfAUaoeTUnQX1Sc4CEgpzA/63dsBQevjmMC6GHdKHiQP1dHIl7qCU9+LTcEp8Md9n
9KxFGSmIycEh+6BH9YBbop9Flw2xwfeu7/J14iznGmWtKgUvKDBnBnhvISy04rqohigK93V11LH2
IhUhDiUglNgdpAZnvbq/1AvG4lb1HDJ/olO/NgbAsJTXtG5DznDJyANN2a3NetHLazfQf4uH+haG
7wBB+w0VUMs26n+16fpQTXicDlTXP4UZwwmQzUtAw5TxzqMWV4pcBKiZgcTuXQRHFuoJ7ieuf9yt
9NiRpn1xmCWfQICiE2cNWpidKEkgxrgVAAVmdSqUT+elq9im2KfB1pgjOp1/OsvTC3G/EPZ4cDq4
619MznRbvC7dfeRUfsVZM5anSK07ngXmmCpwslGvWVSUmswUljBZEX2oYPAT75wNmVk3bp3FE67e
fm5KB7Zk2dtb56y9XrRtExfSKG8ErA1ZUGdQ3fGH74zh+c+LnHw2PspfYZyqoOfBcWeUWkVt5CES
goApdI2a2rchx+SuuWw4uKZwXBaDzbLJJU1/XVriftknY+/824oDXNVPLtzK4KU7zYNURIpQIAQB
PC9J/czNZ//drUEoqSUaqMwyf2evIaScylMXPWGM/VMclXtNs5SEQxBbYqek62a9EmdEHnFX3zZn
sDyYqCoI/9PfGRZZO1DUVKqa8WcMkyewyzjto6RekUThJqegAfaFtm4lEiwIcnvBdwWbcq1b7U0g
IJjX+xffU7MKlz3qJ/DotB3JsQwYCw72LEaIzDr517sv99/tbLvpZLmjfWsfFvDVL4CkTE5HYqFy
1cBXU9hNAklNF46ClGINXKsBpkPjyv/eqzSERfmipfdO2NCFZfrV68537SbbJOKPZKhlhZlVG/Lq
e9H1Dw0a7ze1VxV/QZ4ECJgvbZhIfhf9BAoUeVUq/sIgAWN5F+OKVRe+8uletOxQQ+4I+mNwTYW1
AJgumG49LRy9923sBEzm4YqJuFwBX1YoxrfFOJlmBrnsE5ozCNVHvErW0YZZX+wy4NMh3wWUC+bf
iHuP5bmRrTudM8AotdaDAb2ogN7QYFI0VxbYnIhbOtLsB4OFWnVX58j0jN8Qiitw81YIx2vUBjDe
zmYDxdhZhOdMd4KdO1q5AcuPVaGA1Y7XWKo+r6/VQpJaiHpgWpYq+M0gCX03gUAxwt+H5LtM7PaA
2cydLu4UDsRmLpAaZMQwvRBreRzIbm/S5Tn/snaazjgmSF0Y9G21+5cTy8vgXAhxxf/O5vHm7qM3
6B6dZ0p03j2jEbOWEOzNCJ2hJmTQNDIuezoAZBpWCPHebA2oBpEbmU/oD1iIsbW2etbg2tQj9inl
mapXYGt41lq9fzfHkQ9zhW1TmnhTjfxo+uuenfWLS5PGdFyMiYH1eyzXJNfdcb0psoHfMBWTMUD1
S6liHk22uXEvU3HzL8hAJ66N6KFZOq21b00o/yesOKzO/4gBeVxMHt/+OKAzB2wprcKdyFa5iYpM
6VcdgobAgGV6ITbtGtw9Lm9aFPVbLnO9bV4HGSFaeT57JoX25KgNR1ULijI+tYCdx8ueepFzR4gM
77q2LGl2T6QyCbrO+siHNgfOWVxV223DNmEc2+o/bSFG541p+5+u23accEe3a21scrjN46EPbbOT
A3sZ8GtnvRhhi0su4mFCdaCqqOm/GjNFPh0vADV+xhRx4nehEK72W5oTshcI3s1r7Af8QRNyG96p
TBPYkwRIMHfeyyWAbgpeU+FLtH7mb3Mr3/O58lAjojGi+ydRinlx8NnqeAh0AzZgRN2AUQI5OTHf
KlUm+J/GkFWZouRtzkbn6KT95zXcXIv6Wtq6OdB0DjrHxnBIODGe8+2eB8hN/6kX+6VsD8cSxnai
LlZAqP3/y+kLymbvPYmSDAVPyKPlZPA5BpCzEOSiovaIFLBZTPAipPLI/3LMN4jyvglARUe1pYS7
la45fMJ5+TTJAxuLC3YzWchZrPghc3k4d8uV7dQk1NX1t+Opwmla49zSrSS3vpbZhWigTbY2JB9j
1gWO3WWL6kpHdCr6o33SN3nhG1oI8Mb1EXiwK6mfsRoL49YPOI9/3potBFlmQczA6CrWN98cuReW
+fvxdxVXjLMnH7vfJcy9y1qXxP240Bk4Zt9IRCOeUNHhyeFraUMnMl2yJKDL6umXwBp73B5RmZxk
tMcbb8/Tc4+jxXXGrRSO2HxOB7diSLyXIqKXi4MYGCJ09LjDx9wKf5UZpH/hC61Xrhi8HIZmN93v
dPPRN6EM+ZNrrwarAqKZ4HkZSwwrM7iR68BZsGbp6qb+abd/usLvsPawRPt2oOoicwQJm8exdAfQ
2Uv/Dp46By5vs57lB0V2aTJmU8uzDi2WxUoNCxunAY1dQY0HB44YkplN5fm8dYAzG8vYWLiaURsm
bmW1jLPAGBGwVFOt6NCDiQliNSyKlg4L0eda97kQ1JL8coXnrZoRF70v4xb+FFdDO0wB4rCrI8zw
t3ZGPsT1swS3FVoQ9C1v9gRiCeVkGvMr4oLpnYKl6DCmzBLC7aX3CWHfpDG0Au7kcajkYW37dS23
s+tyAPvQ5vRGH6aM8h/UWzn0hmEk8hUN1lg0kaaGGuJ3236czGzsCgbY9KpO471/ZwsfJ668rBv8
vUffO5O5Kf36UPEVl+now+XdNXpLUfN4qMu9mxfYMupTqkT3S7vQ9wlbaCOmbDWaJVvD8vfsRixX
vHj1qQAqUUJnc63BWAu24XFYkH2NIYkBSeArMTOg3M9vxYYMK1YoqEypkLBtPHDvdDdXwKs1CoJR
X7/+sLco7s7CQkozpX7fUPaFym64qbAcaroXLxKuknXcpV+OuXc07gjODrqiqMSNCw9Yf7rdMeSJ
aZBLFFafC4lzbNMXoaIJexFtuwx/CLU+vB0f9ICxT4ZvcH8lDjalnFlV9mRRzC4COSskQO2BSns0
hT/+VH/4/bYetsAbVfC61aaNB1nNf1gdut7EuHWX9JEX91NXoXVrYf5aZZ8uc8ZlfTxR5UEZ5Aln
f0T4QFjQP47V3cn9sADm6ggmrYFsOqQBlK8F4iFnlz5Prl6h/lsB58pqs4vevSQk6jYPry/mhnI2
WIvoxr+foWBo0vZO8EgK2WRlX7Qv+Wc1gRrYPuL5odmrt3RtmwOgNEv4ToDtcSOkPgFffhKBfGUV
wPRh+nJ2+DyKAXMNEScb8Wrra8eKSP2vJPy8iARCSFql1yALbyQuG01dce9E/8FwM8e+fjWlfiMD
y7qG+2eriFvojWiXQIcwndJOeA2jJeFreEn28ClDnSGn8hNy+7i3Zn1R9tuFounO1xDeKjuH/LqT
w5bmoKCBsfIcXSFqpj8/beJ8188DU+kBpy3nh0GcWQiRlFsFl/NpbHGPc2BVEND2/GQdMdvHuwbW
+mj051NqOiL8Watv42a3YBszbzolkTpkm+GmUmjaRbHjE58/ENzNQ81KkvthK/itL9YEYHbohXah
fcsihJKat4K8WFntDAU9i468BGwpcR0I8CMDiCR8j9ez6ZZG4nCANT6mzri7Lk5F3JxXs+DuwPDq
cA5+WRojeDtXe5x0qScYukeWd/rdYGtQ9fdXGKkhz2v+hLKcHZaiASXOxxDFEd00R1fCLmdJnAZX
Idck67dAxE5NIasdqVFnmvPJ8Z3xWuLFjvmc7I5EdQKsZDwzqSWvQdglXMqdKSf6nSzrBpoMtRU+
Prc7gGuYvTHfR/3ZTm9sMjvxJeG9paucpk/uTEOdZVocuGdscU8xmWYSjzIIDXAHecpW5x7AzkEV
B0ZMlQzTqaim/TBp9+z7utYccOHf432D9T1dRqtRegEkF5jM0UeJMyPzRqu9L/tTXyFBZr/kiUmi
lNXRsue0EcbHlDkvSxfcpsEMbi+0VzuqIxYbhFdqdSYgwgAwi0PMYN1tBJSj20gh4AGfQDc3uf98
v2SXwbh2Pr+Y1S60HOdS/wfYVY9DETrB5Lf53FUc600rkinqh6TSYbzqcDcCTsHbaHKSefcrd/qr
H8knbcf7rxmI3iefhU3jPMLUzcPDUxwSqi0QQy20BCNLyQqULO7UYACSEez9OVKR2mr94aPPYZJb
CDEkIArdxhkLYRJ+JAwV3Kdl5p1tjDH9ryZUtoA5TQXzwwp2LX7CKy09cSzj1MCdmhxLm7nynIoz
DtHPwTI33wTJ3D+UWfD0kg7yCiqdLAGKodd/iWDtqBdCbrC7SKmGEr7HLLnBj89w6dcB9WiP7ID9
hsfwlj/s1Nepj3rUolkRbnNogG7wPkw15wcG7cC0E4wshij8SVs6oHu/1MyzSRRYL0FTuyKofmVy
LFxqk+aQY9he7iuzQCFDc/TgBrQtakM9XwFm8AS8yxbBp+DD8mmQ6bgDUge93SYr02XlacK6e7nc
MUKh7CCpInYa4NmmWLE54hz1Rx2M70LU5MxZV6cPeH8B6idapYVQqz8g7LlmTmpUtgnRtGAcIXLV
fn+CQy0je4YrdrQj3Bd5UN3zF0UStB7I/mJ1jrLeVZXUBvt/Nl6gbUaDXRk8+0qtvHBYEMfQIqXQ
YVKo8lIRhLRy2xM9eGHOYqZ0wcz85Ll14k6eRdHro6pIvwKgQlxvhgyCfxta860LVHzkiczXgo7e
Spj1YLjLJm1j+hfyY/4uy8DyX9rORvVk31e2CU4dfIf1A2x7Z449lO7N/Dk21UPMTjrHp1MPVrd9
0/1BuULbRzDNwqMQtQz+vB2yJyGPL2Gu0NEeRjDQOU4f465Yr9zAhcQjBDO7SAGi44HYSy0OZSoL
tcfOZR+Yaw+vn/gmsj75j/Zj7kwM4EHtvkf1PSEtHSQq8qiTbUOraLfLycFW5FMz2m7bBMCfWTFo
UuH1tg0ZgSJvUgzWXhrutEow5ZrRnQ49QS4KAUenNXmHvKcc2UZ0t/91wA+u31EdUzPAcJOQkm+W
jsAOXEcn5sMRJL+L6xneGKSwXqOLd8rLCmX08xxpqpUiFlWDr6VskjLFS0tzqwdai9t9OSM8hsv+
/zSnxHZ0XxP+TeUz2v6EPL/KizuxcC6ddIVe8e35ZsGlYMs1qveyJq9ItLFq9ROgSujVBZqFA3cZ
zQ7VmiYeLi44cTKJDyQWjxvkbuT/yaPRe/jh8SYBlGNSGOtXTJXQ1gdBHP5qE8U4yI9sBJdR341m
BllC6wBhyDL+H85HwDzKZ6m8Gmbb4Ae+oI0ovhvza87AXIGFiMzfSrxc45ISe1OfYL1bN7F8rAju
aOZ5ijeOkmFajMvLLCSm/EU4VBDmLUH+X4uStGyqwMMbeUb5YcshOkqS7Aa6awV4KROqkGHNvYqR
6lNLJEw0agNyCBzuVIR/qD9lh0UD+aEsWnB9DT4SZn1EMpU9BBgdIObDXUS5ZY/Ml1b5GPMW50wv
vH8Pd17kUcJYxkCVw1ZZug5xfL/OLSwv1splNeC1ix3usm6qzQMF3BAgIxI684Z3sOwYJC66S+iZ
VA/bHrmSPffkK+FZ6b8XlWresqzPNW/88egeSLaos42mHNnKYPUyWz/YpGFrYLmy3bkXp7suFoOT
D32tK71XO9FRV45bcmNzWUKDqaOAr4EPmgIYdTIY22ecAJSOjNEmW+nQKJUR087x1TmL+9LijS6z
fROQRC6Fko6ZmnhevLuPRq9oxK2OBy5atRJZvopyWrszxSplfplsF+ZbRzl9LEe5cNkY7B0j+mop
oRIjv3Z5aDr4ZWDJASQtlwGT5AxF25wKQowkdq0IFCBay1Y+bTGCmPn1Mi1CICkO74zseL+ygL/D
wn6rd/2k5kUB+13ZrIZO4tIshqEZdODpAEIL7DDhl4zZyr5dLvBYYHma1hZcm1v3eiZwPS84A7kL
WD9P/AK+QqHEGyCI4ZBSuyACifj5C7kddxAwTBVjDNchW2E++SxV1jMU8zVOArCFkwCM0pneunOY
nIh0GNa7CXIrtqylp9CWNKeaZ6BEPmm0HOHE8Fsf49sSgLecVTz92DFkOV9f5L2LZWMat/nGjBXx
80qwwPuJNL7W93QQbV12WtEXJKBks0rSqbeK0Iqvq3j53//MdGP8YMaIjFZWM1auXdwVsntaPVI1
4IzYLACs0x7FdpxVEQtaOXjqBz0453rP8JnK7y9G09x7J5Oly2kxp/EycYtQFgSbxQ0MxKAyGcPB
9XzGv/5VVjD7w3kQAFYuFfoxDQeI1FyqIYUqphex0nat6ANBJrqNP2yL7fylqOaLk0EE4keuGFLx
D36PxbQfAaw37GlQzw1f86d2Xx3g87gppkISD14Mmi/WH70wMHoRgOrZjfQMxE8ET/kL2LUs25Qo
p9QbIxaK6ozxRtGH6prYsUYVontZFM90md03/5Lkj3wy+gzFvMH+GalsRdvEX09INkUSmJ8d2sFB
pvijNq7hTq2kPVuP3CUZ1afLC2CDwM8GV6dmrzmAkFKKnP7olabe3hbsc2WDuucC09FhqGGK+PPh
RNnruwEWiiOjerNUxYrXVmZe8jPHAR4z3FN0rCKVQIOlMBOgCnuFnrf9wTXJ65oKIDkLclo50esp
AmZGCO4y0oSVAi5dLSVCPJYDTompMQyEBnamyNVyAJCiVcIqc7aIpqpX9PAgm9rrT/6OwmN1eB2o
X7eNNPrdsw6Kk1e7ICEyy8O15QCuNakO4u7BEEvP512lmXXnoIwjk0UFDf1bscHUHR6Pd1+J2WRs
W3Wbz5+PX3tDDR8HxQUbvk3xq3ltWrRqxSBLY2UVUDoAe5fc9X/tI6jmWB/EbhnuB8/6RdlnwEAH
m5PyEcoCxUC0K+xMLUbfoYs1dUhS4l6nbVucZQHUM9pKmdKBoCtWwO8hESJNPysR2BwbKAa3Gtzn
fobxUSy+XQQq/MminrM13bwA4WSH3VHp2WWBOQnWnY90neTFc1Dk8mS3B7Rev6s2LQnS/OmcwC+y
TnZ2xo/19/Nzc2QF3x/R4UPJDjW9R16jDPrpeqOyE1XClIjSoQ7Y/wssImCdRn/ycyaStX7vavE2
HEI1/rl7hCvDNTSjAuJtw+6WWdektJ+7qnioMwg4EoO/Cp7a4Ytk4nzApJeuL+n6VvO/USHRsHhF
ZJGUzp8pRy/Vp4DOg2TbBWd72v4mNOtMn7aI1pXCVwH1LDrOjXkGwWVx7iJgjtxym4Z2XyTmjS9i
c+3GHpF6Gp6PUTByLy/3sKJ9sr9716CFTumWODGvJww/mQ4/GDBgcjbA8W4UoaQ0MSCCSDUVWI/s
VIM6BfvTMsPJ6GkZ1zIFIoP9elxT11PEx8wjYIkLgj5VMBUEkXFgyLLNInvqDc0hT+/M7n45bzRN
0PZkvlLJmcuzsgb/sFQR1OAfCzY7m03uamMZHkcX34T92or98ciDN+r08w+5zy/WTQ9VvMzoeKLl
guuS5QvDpmTGvhypVa2oUTgjMadAezPgO/uHnZJYm+KvoRXEhMuCYnjykisxrbfKXknhDww6Rp8t
yDqyqp37tW79xyVdcCrC+0Y0pK8UqMYso4CzJSe7B/UAhg5Zc3MvdlKguv62lTc45iF4CK1ohhii
fLYTWKhjjog7Xvx/U9HStLmfyAjkZEBcixb0Y7WOygRrIbHUmvUl1CaeI0d9DZFZcwQW0+6Vnhrd
eZDqedshP8LBrUjogzWDumkXWtfqCBCyFdkl9wR6LW/d8wg2vsWp1I8lTKaFvqjo2UEDWfy6Yi3M
/hD3oE6QXf9l4v71cHF7N0OrpjOP+RidEGyqj9lByZOFKajGflz+cYqLQgYlrHBdblMJGPSY+D0w
F1kp0JSe+co+tRiBPHo6EnMVxuzCtGm9fH+h4kam8ApYZ1SXZHKy22GfAevqdN7a1N4vqbigtzTD
H+/GsWA5In0sXZeMS90uX1CU1FRR7DlYH1jOB7d8jyeAR5b64tfmESSqQpjSZlphGmDzBM9nmTmQ
md9uODAQNJef3qHbmRLD9dR+n8t20h4bizSRoZ3oglA5uk/G0A8d+sgaBJHC8Q+z4f/CKNqk/Irc
c9zuHP4GuclRu7EmH+TIRPExd+uIdFA/01XHhlyxZC/plLK8tlTblwZ8PnjnwiNC6rmgEALqHODR
ACprVdMOhOnbyYxS0ojWZLrdoWCzisnQvr1fFABi0TAx6yEOcNyAj5njGRR29+Ptrc8EqGZNiiPU
J5HpRhDEcXS1oKRB58Et8lHUlI8vQlauCSWsp/SjTfU3iwVDBSNbFtOl1XJ32dzg4nqhGvPUUEld
vK1X5i5oOugbd8tTcSZl7DYLA+XM0c8NTkJZkEocwPAkav/J2xs1LHn1COdVYcdz2ZJOPJxyqH4e
XpUNYNGHvrFPB8NxfTOQCbzAZcL8ZL7v85OQcOLUagJ/RN8bft6KnbLs5ErSwxMnvV9nrPm7eWtK
/6d+fVmDFdJOZvwpRNVI3C2cGTJ9sPwPTDpSKg2SsFM5Na3oiYrggaYCDlH/cLNAK3hiqdJGt1lM
DX/LEuobizwlWtd4oIT+rk9za+dY1lL8BSgCXwUMTzlPI+uYlDScWr4er/caifLfxrZHMVyLnr0s
je7+Gk8jzdKUqVeIzVJCJjeFaRy00YXkyF+PNgQIDcSa+rcwZaeqoJMeoC6O3ruMiKYIMcMl5Dqs
6bV7ei6dD7ZFFZjmWWFngvj0dDmAvOLNg5AoMgwXq87LgQLYMIIu5WsOlUvTZivl+FTd4tmIIlMt
Lax4qvw/91m2kCvnnhG6V08qvVAeNClciuk14eYXI1//r2R4if/b7jV27cgPHCl3tRfbTWpRVo8v
XOOC4BeE97esYLNZw4u51IU74h0/DywQZQiFRh5s1WZA3z3zHITGE4UuUQPazLLqd5BSHm5N8sKh
gormnu8L853Q3CKi6br+8Pz2VQ0x/KAWcImx7x6bIls+DylAV38vDd6R210IPmnMtjYYu1k36iP7
gxsncCnAnnIFHr9SjNdClSD9vc7wlYT/1sCnVh2+eQSUm+Yx602PhnCI3uvB5jUPfQA2TPlBHukO
pFyOokp8H9Pz2Hu4Jt1wRM0XeRPJFla9AWAe0chRw6j77AjsElfXypt0L2OwYHfRkhChHCC7ojPm
BK4U5bIdfU18Q6ZOz4DrnJ2JfTTJEy7UVFyHS24/uSjTZohV7pUqCbM0+Ux5rlcgWdgItijTqfXF
E/AXbx8B+wuuCVZnIzmWCgL8cLVNgX+EN2A0elGQQP63u9BDKj+WBbW+CBQqVgrohImi4/cwFNO6
O6toyJORM2b2tUwsGSplUWfT7XNBqxdxqpYtV4rX3eDSkHUzZC9w6Vcf48ErlCqdNo3k9Zq+poA8
QpgyvHJCBUWkMIJ0OGWNVkWFUbh0gqHsJ5UQrqThkoqFFAwRh71VrLeOMoQ59ptubsos+oL3l+ZZ
UEYahtZ9sbDrUhTV5vLYmP+eEuSUq190dqXexKssW8ra8ymD0ZRLkDU93HLJz7fGvs54DscUqDgK
pvVpvQsmoKzHJnuW34xnUVGLZ0z7I1X3+NHe6x3ScrHElx4mSdjbI6/+pO5O0GwbdPggquQA3AKD
Qqaelzx4XRcHAyHPGg18bOsRM7VkHgl3CD6sBZiWl5Apm2wXecyR/vLOYyyUp/EXBAK2+CLtgIp2
Qv0ZcG8Mwq71VqiQWgVRIDuTbdXZ5smdDr15BN04SEed6+ul5+chIur2vmDtNdyYTFM6Vz6H4CoA
SsjuAyjy9Jz53CktKnpnBW/BQDnnwZ+KMJp6aKRZWAjfqI2sA8sddmyf7J7avCq+fFj0xhLIoIK6
yCBAnVCH6wEfFTyMHxO5K2LntZRpu37hfnvnQ/0bZ21nCVNmbOtvS4Qidhua1ZOB0d3mf0nCZAZY
cuU/wclDUbP2eI73CR27l6LHBaJ93+MOS6WBk9HehsjfME0NMIfoJRy0M0wckCdJ7Yc6DgQVEHmd
Rx1BRpu94stySmcllTOACI1RTToOF5Leo6wz2Dx58zusxp3xdGmsI1f0fhmOu6nliR6n7yIx6Uf5
/Wx4ftCKUahYFvlm7QKNU4pAx37MFb8Jje/6deGxfT6iZoMIms1raS7mYHlmMsGV7juD5BUmGP3L
x9wHFHZ8U2pB9hyxDU09s8ii0WXSFiCmvRpfp66MJdL1bF2QsMc7iG3yPCeVn+ddtuYpcS5oaaIi
YQcGjV7eHm0lRvdkQH2mZWCEr/u/p+KBhEkdDmn8WshVSLzl7ml2KPs3FWUgfQY9bmYUHQ7KGTml
bwl6EyexLY60PZO29LhoQxP12qeOeuds6UuB2r0Ba/RH19iAs7xUCPGfIeZYb1E+KkgXXYr0cCMB
HClRn75Zt3jcGg/ryWcxprMGIZhch2MAc4pXejd94B4Je4tsD1Wn45T/q42hQxO6Hl3eEkjxsmbs
CadviTHMhRPnQy4B5eXBZbBYmz8wV6axLY+Cnsh+xvK+D5hIzspuM44EoLqlNkNFUT3LQ8ug1Pv2
mAd7cqPox7F/px35y+jsn7PGD5mRvN/3Pz0tPUnYa3zlF3EbLVSC94ddA0X7VU2BAezY/Ky+IhCY
f4mUyHk6Jl0s6yruMoQGW3xL8Hse1uNB/D7H4F/XMrJ/h1smIVb5LCEoSI8HpXTmGn7nmGbmxSFH
oh3mm+3xkmgqWxcF17m0LFdAI2WJoOnDvrS2um+UWKv/XgIf8El/5kfLsPINDF/G3afXZudpyenJ
ZUWBgKz2vKD9dYNR9s+WbYIY4v1rBQdiEWbmhXN6BZZuX7ZrtbZ8ywCyP7jHhiKjGH5vANIuTcaJ
HTPB/ZnsSnonhw/2DBQwhl2fdJKhqS7PeRQ1vSZui/0suyTpwqM1r+FvDI0gymW8L6C2ZCym4NGa
v9Abp3WyOC9kHUQuakpNAYCM3T8N9Hc04DOcqARA4/qdF6LTVIS7dGE0y4jZeHkFQHhnx7G8X9+6
B/0efj8DyycpBsHQnmY6Y3WC/ALL9upmapMcQITx5mXzWs8pnbKswMJ5CAHD0UT+H528DicKaMUc
Aeqjbj3OERd0REycMx6QT3KugUTXvipGnD0mzTIvZbsvzxQKJpHntvSwYA3MRod0Lbfp0/yIr8Uj
1t8TYYxaYrmk5AMquQIujg0l7dma0wjEjXkatmLgCdOPA32T6GHZYTBDA7GX4gCyWIYzNdbb3Jyx
2SGGJhLKL+TdZsTkrPq3WQLU9AO6Q8rgCwBe+gNPEyIa+UkQoOT/i5hX+myqchEraKW/Q4lDt/Kr
3j0UQHyDLBZ+WR347E7yuMRWahexpDd3pqUFf08Ec8ydNRm/zZzMeJG71oUU+auc2G6Q/fVydH88
PKPA3s+n3MekdfFRNg/Y9HcEfTi77IWhXhcl7uY40GZMe4VhPMH1kyvun3hgwyO9GUpiBO/lBD9u
Ip9TV7hyrLwQZH/7tvK2rMasprj7qSe1NJ9/Wk/UqlFz7olY7BvIglGq4WV8ENdeAo4VmktmD8a5
kcbxAMQQviNYS/toR0hoYtm1x3m4GFXkvNemAXeMWENuWAjRVN5SyMC1WeIIfBsw7lFKvVRIrE3b
5Q0zr6nk2sPU1TMHSf/YZqAJ8PP0JU63gODgOXsRna67DRGyufBBNlzyt23GkBlRZQ06vZbiNL0O
J2hWgqcmk+WcbG99GPhXqbcjm/b3uS5rora1BOrlcGlThq7lGaOW25iVPfDxkHUx1Ne1wwgz32St
oC2aygaEdRTOWJMIgz//PgFe491iU9F5p29Q0Q5hJg57L3/SfE/ngtOYqosEz6c2iYOUPKzM+S+i
fyxg45MTUhvnV/mIcg2ksX08VReom6s8nDZHgVrcWkFdf5drNKI4BH1OI0bvJKtGBPD4L8vNXngA
yM5faLqBFmcgz8JPgv/kgCxglutT+h16SIAHW3No7vZMwfiXG3IN+Jw7/ySwW6ZuVOVXNdiEox+Q
KPGBUDOT05mxUt1OTTb0EbI+xxEFMdsNGZVkkSvqU7WJkboqhlzqG+lD+LqjjdenzRA80L1ZOeDX
PAjGIMlFPA1mZxkCRFyzzcWJ+ZKlzWpMCf+3PZZblWWSSqjOblxrxueIV3qC2vfGLvwo/clXdr9z
UCZbelG1zqbaYSS/i2fHIAdmMu9UZS+3ffU/r3NycQx60zFmaDm0xb9f1mTZtlwUqty9uOMk1q7N
SCtbXDJYpRnS2ssXtaklehULZBGjHrrWHvhYPgyrthLVHCGboGBLM0pJirbOfI4u7AXAp4CloMIY
Tr4by7MHWgTR0ccsGxKaduXig+tsUy27C7yCZC/8OSUDkTBHLCrhBCpu3G0r/r9EkoSYjJUqFav1
PIOgY5Pe5EETLtFSvTnJ567zrsxhvydBbd27UCEOpOvD0FzgAAt8bPb62ZYdhD6GTdf23Qhfmz1s
1R7Ceu50onX39rp4vFpp/VDPteBzM0zE10Uk7KFroY7RMCwBWbVWZyPn7l5xaAfiNNXsz2eN5foM
eyvhJM2kLyxdPcTm7nka6w0rbLN4LA16a1jHhqU8VUg/iZzLU3ZiIRroKI2Zi4GG39a91raN+72H
b8HAnqfAThz7bMY++r6NX47pmf0VjRGqi8p+4RBnwETTHIMNmjkka95nLg29FOWvqW7+lEMAD0YX
d827tX3znnuvsypQPoJoZcRSpmkbxCJvcvhdSqMkn/rMpNDhtY+YDXsiQu7bbwSCYN0ldmmuyi3E
RAthZ5tCAjA0E9b3uwm7SPdrNOfkHDfVK1zpFM9cCaMhRBlW3VFlJkvKo82w9+VKxhDwm2Nun6/H
uP4CJ8MmlleokYQYmaXHaO1YhW4/QWqItl3dG9LsEltXF/MNBtRVsC8uorIR85nhG5p9eHINjgU+
jodtirYqcgO1kVzmzt9Q0CrPVa9sHePjKuHW9eeaDlrkZznqfrpTZLh/JNyFzwYjXIFFAIVh7W1E
h+hScVi2tFWNjDh3PK2wQgMOmLJvjnNWWoVHSa6QuYIsMiNfecn0bAfyQAlcyjrQJ8ZuWKuTiML2
QNC6IKEbTYgDZUgHKPzvDXE6fi7c30B5PZi4Wf6ZGwvoYhgrHZOxxM1vCLmHW2rXUKRoFhHyhR8X
xp9txgkn0XwB/4ZI84Hxkd/ZdORdUZ0zylmpgUCmgb+m8MIFz62VGEBeoXLE1J40FS33qjFh41BE
i8FTF8/GgnaRtFAOo57jMF/JU0jGBKQnk9hAZX9SJJKy4l8GDj+qbbu2RDr4/Y66kh2jhu/rpsQY
mLS55GhRqWZQyjVac64NkuvMrxYLbJ3qUNCVU+VT76dT/zeWTssYvmusNHgpYSJNwImaRwudiNF5
6PK0fCp0vrl3f3IPmFUvng3A/PKd1UvgIiPFPyllzF3XKdMRH3oOnJLBx3eOrv65WWffnwf87ILm
OHDT46WTqxSwd0Qn2tm/rQV3ab56/LL/N7s7yTjPDeyjevqyUB2veYa96hyXjl28lN66YMdjJUQA
i0knmgaKPrjOe8mOrsTSMIj5Wzwd7DGhFOX0MBtwyJSMHk45vF/8yMZtM3a5fMHgdOfVUvUAMHzI
sE0o98oVNXuKkS6eXKkn3feMWN16ykOyisbCVjH4679aV2Gn8TExJAmf7Lju67iSU/p9M3voD3hx
ePtZRXC2zCBd/vSxYANyWQS9orLB3ymqmHh+6duVG0tSI2g9lxlUcaYyaKuPW8p3JOYIdkkWhwiU
YO1IGus09vH6FuWNw1I3Q8vmgMhExO0hbk9nGKRmCX68sOks9a+wmhvwQ3XNMSbCiODR92c/zfZ3
u7+ZpGagnCcRhUmx08u6Ie8itasbEgQfnhHQycsP8kuKlXXlXQU8BiVDu4jBxCG+PhrjpnMBDpmT
fwItg6GMdhh2NsN/o+JvYO6iq2j0ArSb4QoH3PL+vybd39fH6aXUJ/sHEQI3UnxxnKQiYvcDQxbY
g/N2K8T+3QiImOF1J+qDgGirAuw5iwPjo94SixQNLhEkWq/nazb0adPkSS9uHYH9UJ006dtlDWA4
n8AGxVL0kfmZKcjvb/U8G0w02haSQ3hUeoQLmcKtq2M+eKeGvbUW2rxI1YB1c4bJjt/P64//aNnp
4vlW3s4zRhTSiLsF1GsqhyGj/RpjYEQQqXagVx12J7oEKXv2d155erg8qMk/n3XeRjq98vCvNTlE
CLppxezyJV/h9srToJ3wD7TSaZXZx+TepFksQl0nUuRMj304aHfDYr/7NZGNHCJJPCgQTP03j+CL
XhhPJ5N4gcM9RL2KofR6Hi2dGSAd5GUM3xmDDgyBXwX2JPSnX+6JwJL6JB9JSkrGRVI2xGwbK8Gd
YdR6EB9JrsMNTnpWCm0yfB8KlNOofOGlomnAHGs8RpwFFgbXhaiel548WVD6rI1hgv564k+DjIhU
iDD0+ZejCwO+aKpihl/60kHMhw02Y0gTziwOoIMRELyXLSWXVXI3GoroL2JZ++ab/oGaJ8MihsU5
r3afqp5FUu7msEVXqrwEyPpE+1Ae2zcIuCr6SAabUOireXWl/5qWC53Qnqi/wa97qndIJxIjzZXc
siFbIyiP3CO/u/iynz2djgELecpdhvz/VcMJhojRBIpmjWAaEdPHtbTuxSulCK0QGuDezqElqJiX
phvoPjqEiKVMUsUroBrwT7v6j/xxPnzTjdUrJYNnasBhr0JemSrs41af6g58NA2q76ZN+SZ7lnGP
QobyEBfgmyPOt6FE4+7HVEYXCPrYrFE2RblD19iW/qf61a2hz+0KHKjQiK88i1+kSV32fIzKIo3u
5m7eEhs4LE+kOAAj2bzHo6DHF6rsBliWcGFaBxPEUCRciigX+13nizH0LX6bsj55ndMKXOZToZyv
40rwuLZuAX/wQ4YCO7iLE0LHMhQMRGijEQXdF/T44DG8w54bwZiWBZVumw7hCxhHUY8qBlr3NZ7R
G6gogBdfSLgdRJ5VoUmPY3ZUDHOkvrr9LCYFj17n6rieDQMMZPsgC/QhfsLndLvEgZNWuGe9gsRr
+iPxAFTi4bvadO7Vfo++Q+ckLRMZht7KCJTbw2Jwg8Mk8IMAbvL/QMQ0vO4ix2vNmchzmqF1BXLw
G4h0sh9UL286Rj36nmsVm/o5FJ6ucpKXagcgpE6/EU5Kge1UaX8L1xv0YMz3rbQKp9TTAfWdiQNn
1Bo357S1Sku8OtC1luAEx4aliwHJgRyJMeuAI61R3K0X4gXfr2FpWUIPuUzEL7KzLExhTAuBbze5
QNKDqG3vWZXXM21NC37M/K5hp2qYgdGdeOqbe5PwN12hCBnQ8PVfx15dQXpJd3LDNUCR6pVpixPY
2GmYvt1KvlDzWq+VgQibd6mUj709s3byhursYcytAhq980uvI/6IuTML2SimuFjsoRA+aqDD0o5s
C+k4Pt7ZhZLn5ccePFWxX8ZwSS+BWPe3UqWnj+qblWREtAqLbbnz+LliI6GFo8/PAG5v0JL4qjqm
Vn9nmkV0PtYtBWYRq2Diw/e2pbZvQXMDDTHc/8cOTJOcymKZIDheCzzqhr+ieh/B+/79+zBZnUEX
+QdrrTICCusOq/dQjin1j5QL4L4HBvf5vqZoM+hyiO/pj3GRLNDb6RYnXKwifFxaLYgrVCyCTnFn
EyO4MLs2A18XF1En2ywYRKzaG0wQWOKO9+wuADHbZkZU8Ceuq+PqfCWUmC9lqR/JYD0WdwpKN2v/
1Nt1CoXNzcpcHzMFD+epyIVtf7qq8rprj13dl7mRBK06Pa75Ws05QWaEM9JXmg+YWZeauw+e47Ay
hNOABXLuddxfIwK7dThAiKkqe++5EkPKIMnqKRrHmVbKe8vlMuwKiROGrbVOpPxzQPkFarh3oJgZ
pu2+IDdyKCMJn6sC/Jgh+ywdF9BMXOz3hOw7qofzmSHh/PVvvm211DTTNkdg7+FB/C/n338nyXE4
CUvPcUzp0c5JSczlydNGC8LVLOZRY2nmJg21kLkOOTuu69LiylT+xJ9DIYfhQ1IteLXDQ/73ofLb
XmYeqHJadewORdzRG/VnKFmhNFMdRyAmHymPEnlNDtiMyVI/e0O4eS0ZUeuRE0QdMX6gI8Hob2ON
a1/Zie5nigYgH1WlDcls55gbk9+RT3Z5KHs0H7l+7Ak9QMsBH00U6m+/QLp5yxcwoaLverd5TwFL
QPcoc/UrwP3ONVAbEpfWDQ2eoibIrSI/+eNgBXqeiDvWHOk4O6WjVGmyerb+/ETzgM4EVpprGqaT
sRFvllI4flXqDN5IY2DnZZKJO+m0bFSe/qy7K0VD1nNKNu8EkUVaDRHaDnYCmysNzrCdVPpJfMxp
S04lkJ9bVRASPPDGQWlwh77RSbCHGBexqVyyzoQuAUTgbivQHP+ss+Xcig5qGdE3i7PJrRhV6zoh
eHsZv6JDpKELSAVrmaZRD52vdZCMjnpXXNv/0HORt0UMLF0lMEspXy5VPHQBgx9y8cOgUjkxvPaL
5EAxHTRXhP8iSYUgPbLWz+hoJQs4zHbkUXQAlVEns0DzT4+5Wewrt/W47iGBnZm0IJwM8QKNu0JA
TaYHIhzwZ/TqPO4FfzNtgP95BRIJgz5tfFpnkFJ4vIKAL1vwlSChL7rVwdtIw8UAJH/iNoCvWZ1R
B5m/UAcHELKReO9OMmBPZMQueFKhalhMyI+mZq1hnWhNpyK5ubpBQdJQ+tYEuTwG2etR+rj+6CRI
shOsOEaOmPcbJO/gkTdv6+ooglHAZYeBRB/tyFPy57/8hnmxdEhfosXmdmPyC0pTj4WG3bXsUOV7
MBbmJT7KETwOr6SGSzb+ZJJorpVxJvngy39fagN3jbDz93la2YlayWGorHahHIJP9fzFoZiguvk4
AEsB4XYc+JgVfsrMuP+Btp3YUPkX4osxCKiIcY/cIBrqvDgOCN2yffj/JLLVFAIVChix1P61DlSt
d551rPTByb8HMCR+MrWMzXSiJcwzVJENNGksBXRyMy6nv1kQ9Uj6W889/8QtYGYa0X8h2aXvDTcN
GoQ32Quo3lv7onj66yLZ9FaMSiug3fr5aTRvha8V/iVa3ueZQIbdkblB0ewr8gpT260G9BNQLcCW
iI+uuKnVkmC6f/FpVWE7AwrRhYZMD5oOX4vHOGfCCCJICKDYmdko/XHATeH7YGbpYKx23vOq+AGS
Xf3au3jiYugQXISBVvecwLFFF1sCj427ydfpA3pgRF0O5JSCUQjnHIORBUoAdUCjZM9logKAedni
8FjbzFegU4XIz07PFr4ll2hMGXlmTTv8fwX44rL07+yRCqTQP1p2ubCPm7iTxcGQP7fIRbpq/Wgj
dnlTJ6ymOy4ngRwxyIj5pLo4zDP12+W+25Rwh0BLCdPi1BG1PvshYWmMWwckkMqhnmJCQ4LTsXnQ
AjVSxQrIJz8s9DbnAAW+xxtWTpLAEUwDu7jn/j7z7OKEEXSE5CdHG2k+WacUTub3BrsKk6STy0ZG
W3zg+ONkkVgRiUuiPF3cJ4cVtQoXEmEfa0a/+BUfbUPThaTaCqRvLwTIkJPbIkhjfp75bqEEL+a7
EzZzjCGS5eJTcTGjAky80XynLMnx/77pdKZOmNLVx8cy5xZwLpVQxCmvTgYjoL8GnSRMAhrMHB3G
oJD6ChWmrGd0PgDrTcs7WdFbDO/xTr4SlMi9lj9JjufmxkMQVxkiooCbJcmA/FyqOJMPkl7u15rZ
BSzYxeyWrFpopdk5Hz868AwgBP4cAUNaVuROU8qxFbt+El9UNBWXxlaS110/xWBbi2l3mLY6XgtR
s9MdZZjOqroOQl6quhBdExXCwQCe+GuP9xVGMrXrNopOj/rcanb2jTK7Hgm9giFDtZ7Hyz1g92UP
J4WYhIKmN/BMJNg8CDZoAxkjbuhNC3Ishcb1GLWFtT6S23m6SyvyhsZkZrDHeVWSrPBK6JoSrVjE
bFMkWkqdHyp+JmAq0VoIYPukx9cktUsggTQuHSKoZAc8yhX1/9EsmMb5LDEJS3RIQlDY2lNloCw+
HRFog/KeIOf06HHPpRZVK+e7lz1IHGWAogDTvoV0pQPeAiMs6zjQpJb8dlqPbX7bE+gbLSjRiUJS
gMD/k9/BjmTf2l7FRAI7S/ZRDAnpmrVfH0ZYolDvFJSNZ3ViQniBvf+37rJqSL00VYF/2TodVdqD
YhkmLGs0DokspFsecwyPEKcWNjRLLlb+U3o/24eX/rrDmsOPB+a7Tlovy0N6vCjj0LVzn9kDD5TP
yao7rMYmZBT/Ne3X1ZIKnlnqp0fba7ulWbY78lleoZbJUrKWywXtzdUkV5yolEhBVTNMvMEgBD4W
o511GUMo7Ly/ENdpFSHh21C1iJixV3Rv/JU7UijCJG9I5coFyom1iP0OmaIR+jhqXZmnPNPijVw9
tKSS/IYILX+aPBhA3Pk1dCWAy+luV3PaVY7/WsLcw9VfKxvFefg9UEJZ4zhybjyHH4dEY9jvkrwJ
nThWDtZQ18xCw/8Pk7XypPRW66LixNtyLJxK/uyvfL5gPmxYrhTqdthmX3cu51Sz4vpjRAWVrkKM
xjosOI7JL8izwISooO5kZTHrT4ZO9F5QC9ndSpd00TuViJGsUewN1b9N2pAiyOhkps7+y1yRYYeJ
g6Jm5rdoIwNHq16VU1v1oGaoQMbTy8QwUsJcD44utn8rIsSf2XOlzX1kuigoCRDs4CCIS5UJKXIQ
w8R1ZtW4qROkm1utSfOQZNQTpvkfrbI5jolma/Sm5WFOJ+X1I0HzTubKjfPzjW6QWrxK5a+EeVAa
a0twzdITn4Sj/VBusT/0EQAMHIjQHM/1WKMpxFZe2X1UjsFHwGNur9iM2PNBvv5xq+0xH6pKH0S3
nxP9yV80suvEgX01wfB7BwKowysfqznBpHqd6cti+vH8ofDEzse1yRHoWwhRjQj3Lh0/31zyTbbh
2jMFBoB9epDgcuQ+PBpy+jJ7cuY3VBb6g6prKlr/JKpiVrURgaMeB3CVia6wvnmAJD2g8urAhpLT
y9mGRCyYx9+GSiOHoEHLIuW9EiGJayuIx5s+FLycS3TWTTW/WFIyLR2psHHaj5K9fmYxh1cTvY9L
EJQiRgKksd8h8whAv148UUs6EVqRyAkF4i1dqsfFkc5Z3bDB8Dl/PRpf3jzMbcSk1BhNioMYohoO
xbm7to9PqVzNpsMMVtCrEzOEUXfpm8FPNRDQk3GiS8ztuiACtTcTOv8W21p4zi2m+t5uX2S93c6r
gTlf+eqvJw+U7Oq8OAen44KbmAjs6auGkVQmdzEwacJbjK5Zx/5y8k0BiJJV0/g6EODVGMmW+Bwj
PVwhpfb9QSIdl85Hr3b6LqpEoFHFRJc5SO+JhA+Zs1RChxnUmePSdUZWJu1LStdaJeW0VteqGaoh
S6JderSU+wcHKg8DBtH5NqPYTmB9JSpFimbKvALSrraWVQ3qPFaY/qqu7K37gKE+AoYEbJi2yr8d
b4bDGu4t5rXzIe63Uy5o0iHnHSqXVHfeWXGvln6lXeAqMdMU/sfbN71815pNNvWWqqHx0rXCPWG/
TNHjxTOHuFGmM0MfqBbOB9VwgZm5c5PJX+XoT6SkreuhAO9zcHzkElNl5/+Xxa/tRxpK0SZIdjHI
MFzcK3mtws40hK9ZtsaQ62THqwQKrgCmpHDmraqxDS2BWK6txRo/KOB5qTPOOjFH2OH7HkbPOSej
zifKcLJSSu9BZeq15JTI3Vtz/o6iDdJW7mb+U+aETIoMR/pVeRM2WV5duMYAzutH6i1SOOfWrk3x
PCZJFHJFxO2WPPhO4U5Ml603UNDUFI2HaxrQTxhaqm9tpixX5cOuC/LpeuKv1jtiDW+rYmIEvd0h
tetCFHgFGPLp0hZkhIBk8ocZNeiRmoh0wMvy/dNlQV1ZL3USj9QiPLDNheXGueYmWa5lY9nOpK2m
eBHXB8JpdSaP3nAvaFPc09LhltqUWT3ezhUllmJ3K3Vefjpr/ciG5uukUkoKwU1n4f7Vy0HXQY+a
aOz0gv2hxQ04i405ET4+rLaAFENtqjZJbaWAPTW0MySAXWfg3hM6TdDYPmH2jApdNunyeZb38msU
iqCZjQ1tdkG5nKrDa6H6yyn1OUb1Bfna3qEmSfh4Z9HkhCV0YVdn9/LVYLvlJMfnpClUevavf5Hj
KT1C7oH3Ly4GzCDZw2gJis1NC148nNQKjm/uLEBc6FM0tS4CnbIWSQ8hFCa428YAagZyOYmJoRfm
f5ZKYX7462qERJdjkXvfQruQqkh/XTz0PXGAW3rfrHL3XoUhDIDGRJLaCbuqwamxAbhzEebHGe8J
ljyl73CwaXDiIKGoRFmrb4YtCAO9ezALNs/M8t2oXyBePZxxquUg3Z7GJkphY3toYWtBv/oBX7Pm
FqQjTzI5ll/jiQsvVaVb+JVU6/X6g9B83pZcxIk6irsKsGJC6HiWUzLvommHk2h5EpRCsWSW7HcA
OC8xVbkltqzYL505PB5CqrQN7tdk8F8Ma8pjujmBl8Q1zQ9puxUnVvU1qrPIYclGXleZAFLkDWbZ
H5hO4vJk3C2GKsMvfem/FBe7kEPPBcp8lAZBtk5r9OjzidZgoaui9OyTboPLQeDrLNDDIFr4/8rX
ivYyjGxgHAUTVJIDijVSuUhjiAmL9ckBBEQp4Jn/SBZfT//jbvlp+ALqbuvUfNgZSo9+bB8vIjQt
/DB/AVa0Ka9fko2MgTbJXt4ZMGpH8n3UIoB6QUl4BhgOEX8PQx8V3e0CIt169Deovh8eYPzAMWdj
X0mT7eUZvMCvz3J/Lzk3/q7CBHxc93MUSlxD4w66noeeze0yOc1VgIjpGxAZTbBgzAzXTNv+46Kw
8l0lfFyDzXQz60/efRjMR/AaV0yfo6tq+ONLr1bqRj00uhEDSkfOuvUM8Ls7D/8YNBfJmAI5Umld
XC6fIQX4GVGzqQg7h64h4zudnzT1FUk+D1e7lHGKnrmAaTGdajPEUmYjNfmHSsx76fcqr5u7gXOs
1Q/8Mee5Tt06gUzJeB1hX3zWqWGt5UnJ2aauuMRi1r9no3X4I/b8rJurLNEEere+SFg5etCLMore
NH3Y/zy+KxVeNc72C/9nvThItOZIOOiZxY014Yb6a/HGrSulN/6/CL43t8KXMPKFBZCNl+z4kNjt
FfVf+jj0xbT1Ij6tBGZGO8vWPZGHIbEszBV0BI4VGhGZME0CMDHbgbtGg39Uz7a52iusYiVsOAMj
U0WXceOuTKmWxNuh4EuCBUyduiahBHSk3jFoYdXn9MbNeWqJjSgwArazkMa0hxtJbvcqW0TkvDjR
Iz7z4F5cCSSrE+1bBTmCB5hkFg+dtiw+lhqQhv84cmB+va3Bc8/Nx2yh9sCKdGTFpRO3eTj+bWOp
XN8MsqtGPZh4d0/I2w3zeqt3yQi+6reBVQheI9TGth74AMpf5QVjgpvFOYOj6v9PUNuv4nNzXfto
cjw3ymIRPdIO1ia8U0A69yelufs7yL2+wlNl9yI31GMBeeKXGkuse1VDMvSSi7koffiv+RQfogrt
vAhbOCdzhpZWYKn35TRfMffSK0H3wrJ8TNMBMMBUAvGDj3jMNyWso7a1+p9CQENfpGN3Fi6D89NM
SfxTX4WP620LhsKwkQ60MF80jlmlvDnBrxsP91yYYMy8D7QwBDy5IO5gDLuC3/AK8dxboY2LvqvG
RwwHzzWytzYHEXmw+0a5Nt+8DoGHU4IRRv6ezKwmaF/2kZL/JnC1kT50tNDjpCVoDut5ZVMiY1N+
voX5ELag82IcK3YytXjLFDWM+O3DEJAjSlBQ5+w5xCyaKlQ2EqPjlthsiwQAatjZMED9MsjZEN97
JH9g1XITv6fjxPFxmgWRmnf65Upm3sVNM3tV7LwViDborF6sEW7C8CnlXc0jnQ/EL5C8jOwRkQCa
3OR36BDfbYP11Zq1o7x/tK9dqJUL56HaqbgQJXYKVE9HDpbdrlivqAcwJBDTLWYDhpJpz7Dsl+Fd
pLFguoMZ/XPD6osy54EUnS5VGoSxONK6gtkdrgMWpzZwLiptvBeniHdlGZ4rRawjOkkzbuhQtrDG
d7a9uZ0jDdpDxCT70gkAJal1hDwzYU/LLYEo8UXQIPAA743oPgGgqtft346cnVLihfskThQujcUZ
H/MjBt+xnNQ9f1DC5eIxbUCSEAd7cHGAuQsAE/6YFCxhi/yTTqs7G5ozZUwQSkXLoGuB3dJdTH/F
nX5zQeeCY1Ad89OoKPWq4WyQKn5LWHpmgGg4N1jzVJg+U73HKqSMEAt+qbd/divnnQC6yUp5MUt/
vsw5g+Ubgpx25Fnl8Do6xe75F24qWzeHyGeeL11esSCbPGy+KH+zeuYjh3G/QI3gpc5pRXLfGRWZ
bKWYgyBgHbeXUN96lx9b0TIAUH8DZZmFOyd84wGiQScvy9rlSqZZ2+SOfD6L7i8wmcl3Gc2BjQsI
0Cs43EHLyGcWNaug0v2Be4Zngu0/mkFugoTjCQwbVhWHAcZRU4gUvAXi2IGSsEe1bNrQ+ZRyL9+s
/ZGPUUzMbqwdYXBC0S6u2CyQ+Qx3aPkRLwmKs2XvV0DwEDQZp1y5DlBWXmH+gMpQNntikgj23Fal
8MKOvzGFzqP2a9W3wa2zefwyBGg/3RP4Hmm3ZPGXJ18oRYUX5gisXaZYiEXvpduvpaIsbgZ71P4W
i/Nl/MW8usei3GEZrN+y+eMFA8zKLC/JJifkKZVjH3/WIHlZ6H44tiuM8NDDB/q6t6UXkfVCtl4V
SlFfF6bgkOLIt/K2urxmu+wojRTutL8eZwQmoMRhW+U+x15TS3JrnLlKeOnCHCELbTh102p9wAYy
tjd+jMFWSzRXPZxG+BHNqYTPVzyFsPCntIdCf3XxJ0lyW5gdOLAzIFdlueh5ePHAYahZSZMyC3lW
bzLx523al34xm4lJvJ37yfs2XmLFYXiinibC/vBjMXVa4QBIaj5y6sPLd8SfE4Vj1efD4UhIfP8S
SZt7u3AcrbbHYHXaVxxaI6qGNG8tNZ1uTlVWWtIKyuAUryxgy2pk5NVmcRoywIrGPB3Wz5HEh7Xa
BJFNEKPeG5a98L80bmwrFYrlp/wMRJh7KajrGm1IqdniyhaS3Sd7E0hL2ThwOyYy2l3fqCWbnL4s
6SnG6MgYl89N8qR+cJ4qJUy329H1JYjbRwMNe6hdg9/yzpJLqDRiEN32N7cLIjzpQ8dphqRHrwE3
nIJWBS99X7oSkHv/lwuxkgrOTqphyH9CtzF0qR3LytZn+hYsysKJSM7Se+Xm7rQkEcIVuGLzJWvP
N8C//dY357lGNYZC1qrg+qjmYaV1Ee2pXr+l1JKk0FbWUVO23rWepCZNK+DDYCXvBKjQhtgxlCXj
p7xoE4pffO7BpIDZtkpaYO6Zj4acQ/3yLLzT9muUxCRzlIiC3Eoj5mhh9nC1i7aEGNZKsIRvnLYB
3kSe9JxUsyV2WiTM7t1fpofmLV5MbRNkINADqXKLF/cnkRBgCE45eXmPCe0waSUD5K8ghRi/WOMq
dL0nkvZ96h4g3QNAzEqpkyoS17i+KUouvcxwJSlzmGB8kanZcOZyOcMcA0AuLEQNkZiSg2wxaYko
gNp2/ionhfJlRGcxU25zdgXlusUtlVEN5QCiu5MclrvnhEMLLZq6+mfG2wp4XbAYn81TqhHfRkcI
7jTh9Qflv3TCLin4qU+f4XhZjZoB2iDL6DOAzadd8xkj2A9mLuwK1qppfpaXJ0B3aOIYVz1ZR+Qu
dGYAps9tW2LYPqbjTfY7y6Oqe/dlPuhsn5Vz/lmEdY0XKNppFzmHNWpodWMmuA8HEUJgMU3NPwGw
/5MpGqpUWuitNncIEbqmQHKsDB1EemIV27vNrbVVrKg2uBeHIc1l6k2SSeSszg+TEjF9aeEbnFqU
2Y3e74NFxZS1r2QKRpfQhegtweU0zxUoYMJXhSz3I9hx5vudep1KjAMwkoPM4bqtF+EpdWxiBVWF
cOZ8xHA0c/bpUwlPn+VMEPjU8t4AOniIwLj3pvU853B84nltbegm2S3x+dVbbKXlhxuGVsmKjS3i
9bwirr2Z7OHkYZZambfx6ZFjCL8jNF18aJ7NbCFUiT0cWz7H+S9MoTa1pfnBrVHon1bKEo1rZE+L
4HbEwERia+zfbxhr31RCLlQdZwXrvYTQ+UfqsDV7vDCjpxggkSWVXj+HVCw6G2+9/o5tLGPSW/PV
hz0GJ4zq7iatU6qvCoiQZaI0bQwzphcdgyhUYVOM5E3l7L8qL/nl4xES3fOsWf0EgCzeHmL91W3C
dNhZBHbJVjnckTDg+PEFCri7y+Z1ygMKNtVHsSDUR7RWsfcmfFR2f7TxEjrzL5FNvbmV/FknnPzK
bHp/giR8wZvokmRbqSNMePUj5Sb4DalK+pKe+b7J6Drrp+j9CvbPEuJxmdetwIl9eqZvaOeZ+t6R
fyRO75bQOiRLiKKUWjoUc1p1EE2N+Hix3N5g5EO/2IWACEEZwltoroAIlRXJGuvpMgMfHMWQbBJQ
5tzmRoPeVDG5+8omnr1Kxuc9L56A26lehS/0FSs1JXUh1c3HCnKt2jQDcxoROpvkQMh1ePseACR2
0sgM+zXf1n8u2nmu0YY9KH2dbZIjIuEdKKsma3PKpGxa3VYHp7VYlXfzqtu9RqXBoFE0p1WOdEvs
V3YDFwWMaxO/6umy9Rr2oBaDeWDG0bxnOly/4iWP7SR0wIaYpwY5XhLPvhWpB7BchgH30ZRvCgoI
ewERISGvQNIGbkiQDKygOJjDpLKPIj/wOhdO1GqpHVJHq9Id7TNjXjOiKViWxYDIQ1r/CoEHjbLT
nJ2+E4tvTWg6K/4Syqt+LDvkIAKE0A+6WdG7AFSQqVdWiSxR2by3MN4o1A/smw0AaXYxUt39eXsB
Y3NIEwtK9l/WSVjiY+DmaFfTaw6TXAt/eoueWDPWiYVV8RSmU2q7AWGQH50iU6NkdlbHgKHpZuFE
i5u3geXGgrD3H7YLAXPKJlX24A+VMHNWEXVQzOT0UbpsdLx3A+iUmbRCewnH5yKuG2GtxvLO00YU
/whKwZqd9sLJcOOvkeNQcXSDo8Mt+8a1tRi2p9wOxLG+Fx8hUJG+ZON6YG/BI9qPjX7dym3Nqtj4
drN6dmm8GlqvTxzSx0KWh5j3cQG/t7MDn5/2gFhgUEmQ6TxiDUoBFaFvG1YfwR6e8ZdRpFtNvohJ
jCtWgYTL2K/SVjcyUCfsvdgEViGcBOgc4QdhQH90Tg7kfgQjy7M7q5x20Ks4O0CcMzGWA/7WCGEs
OtgYFM1xlLbWQfclmu2iMKP24JteNNVLqotPXkhSloSOk56BlFF1LBmkt5dX/0sKONjaYaaLpMWU
eC6ehC+qbi5WItQoIGqyMoP4adZ9Z6fF94KzNI0Sz1kwQwy1rr/fWQh1uJMXhT8EZrYVmHtp04sy
U8qKe1ZyKa5N99YQWuWh0fFEOLtXosXtOuHPaFDjhkH+CURm6iH3dg2jZ+/3matlFu2TvLtf0hfY
tSNU7ffVARxEpYl31GgbFcWXIqJxzEHmabF+6rOtUOueeoOG2vGIkWsGqUUAxvrBmyN6dpFsR8Hh
zFhuGfpOOtnYPqEuWnB6TKg+y0Bp4r+n0kZoZ8MnLXl/gnBf9tuh/rQbpFBa4XN0qjTOsERp5WmY
LdE2+Vqf5Oa2fQ9nTBYJfaGcyieFrBXlJApzidqSLvwFKAbYEAeUOvU7pkgrkLvHwhPflEzqwnhY
MpNw8CQepT9+7hncoNknKtUXL18bPfwOml7khrMzjvSEzr3uKay0I9jpfJsCkjlZ2jTGAZNMIHSj
ELk4mX36/VNkpO5YRLAEa+UpdYpQDq1/0CBNg1uysFHm6Hn1kNF25iB5VJOhLie9VzVihALmUjub
YwZeUBAos8oYp3OTbBjRLpmD5KF5/T+6nTepTAfiPqL50q2klo22zfbmBOhYi3NwbBTAvaDdaUQi
AyQjz4qa9z40Qrj7QPQLjBVJiiDecopIKDi9rotcdM4nulb/GFF+lZqGgj5VZdq2S4gIDgCA14J+
d0fiOdkRd7ZbOPFIuXgae+YxDkZjnWS3jWhHt6RUXFGEyEfqsgm1FwSkAjbCzDDqRg7tnFmhxA3e
8/Sms//cONns9tfs5iUQWW7nlhMuXPjM34ZqNc/uzW4JSJG47slGJmAlhoP5xiqE/oqQp7zg/vDo
3mwbrYG1R6cXgq2uU77hh0Izr5hm9T9ekIGDJ60b0P8YnYlAM1LKurGBEOu88iXasMwmENoqI/rI
uWZs2y1KjTJdKil/WXTi4NtrJVl0nL7fdZbjcPyfu2l2wZWCnh4yERc/ss+43XpvxmFVaPqEH7qL
h5B3pBcpljnr3zZ11H8nyNAyrt347lte1QasxyBfMJnaO6VbqkppKJR5Egpk3qjm0eXBy/Qfydgl
Av27D//8sCdT/Ska04NnBqlO+LEUVgPct97yx5fR6aUEXFgJS0ecgZyM6QTIDp+CZdHe3ks2B2S5
a/AYt9PYVCvg3p6BtgzO7V8LnDh/kK2Gbv+5Pla+WB86CGLxDeq7TPaeKg8eoY4BmEjEqrWJ21aM
9n8UNj0fdfyycDhrCcmX8vx0k51bUZCZE7CdXkVF19m89Tk+INbmq3hvTf13mZXMQz5yVv5gBcP2
PDxz4bLmayC/ik/iApxE8he8g+o+xujV/U6uAO4YCJsXuBlEXEhQ/HszO99o3RRLwSmSc8VTO6z4
xbQHaK3xqIG5PxEXWjV7JvDWFhUpNyrV7EU6Roe35YJ1Vh0oGgT7dIlKydhU82Y7meLaknVXHvGR
gLJlrEL+eQmgAN9jBHkohQqnetxjvseEMpnt/ru2EcYmynxyMNBeNTSyQ0CRUq1jKUy7dnpEoOU5
5Eddvoj5NJfwIyAo6/+mNW5aPdJcWqQQuDy1qkrXEEiagKsCAvWWiAALa4563Jvg9pjRUTjXsC8a
AqyY2mOzsjvL1LWjpBbbb0tUqpD1ku3nXY89LdzlQcarzG62eN4/qFk4UWE1/NgVQOVsXeLAtv1k
uIMXdY8OctA9PwinuLlDkAH4PWZIfKO4aT2bjyVXTfC35n8LDZJFQ5EBiOWosdEr3bXKBtLBw5fC
JCSHbO8vaE0VzprDmKxNOhMjKiaoCO4qXhs6oUGf5R+5c6SfTIyMk+KtOub7xb3QrV4x53zBfF1F
S7JNbfCi1HQJkRofA4gOj8qANrxgQN8Pj4bf2iefx+AY7yJlCOLS6+gfoFehx4ObP+BKOPiA8Fn8
GaLE8Q/bSDzSsknu4K3uuoO4HAQxvTiK169D3pGOtvb/lg8V8H07FZ6uATX7xVlEfjLn+7pBjEcD
ijlyl26YnUu53Kyh463QIdoid2Em7OZmK59dq7bZG66m9oMJzb/OQBUCy6Lyq3EbLxleRpfrlGl+
TlD8L4FE+eFPBRplfRCXgMpQFvPtWcUekIs13XKgO9hXBmuOEzJJthgXdE+78j58Ngo1eM7KT4Ol
AUBRpDIlBHZ75ni2HbJ+nKc6CFNTRSrfN5kQsv20M42e5/kllBCc3k2H9gJbPK8UuFnYSnKXxWX5
tpao3SRX5IOp9XuXgn7guUAg5i/x8h5qyutQmLiVnQ+6Kdmhgq/EGUbcIWORw4eOC2a0eg9gED0s
LwhIXm6uY8t2zEQpS7fdK0LnugVuoDJH+4D9fdd8/jl3we85nYiWVjSgXkUbqy3WF0oae8rphPP6
Qvx6DOgk1rwZINfjo3hfOktlpzAI1c3xg/aHsu96qWt1Dwphet0k/DQJlPsKsYR6JhMkCaGMHWUU
bpyxNzTHPSJR3kbhX64Kq4jz+1zb+QTy/mWxLmAs4OhWnW61Ij9C62h4GbfGLFqhN8YAA+LGMcYG
MsEDy4kNGI9DfRcp2eQ6N3wL6SX+bCNoSpk5eu+9/oLSnt0yWvTGBlVQXOvZ09VWeUc4xgDbJHZ/
Shrni5vsQys9hy1mLDdOqPcMlXpIKNuCT1ZtAeJ/7QqrUBkHPGwYVlkYlz6qWCOwsqPkFhORmQts
L+gpEFhHf0SFhyJMq8Ene6ZNqgm9KzQZZ4dlYpcwwe1tRNZY7D2gBjtCEYpg3R0KTc+TbWlpiXfE
JHCCKR3Kfkxa40jHjGbVP011DgYaskSGicxw8yM8SWJnasx1VTU0SWebvrQGRcOe35MLu+zZT1Uy
A3PMul1eDlj2rr8Tefsy3/oXtVVcBSd3rSLIqHjnCCT4TaYtaqPCdi6lW3U61vQi6uf13lbS72Ej
HAuaH05Q9eTONONGvAeSxkgYmo9Ll0tqi7aHalhBpD+0crIaqHCpi0vYBl9yZXcnDx8uaqJ9LOLb
rtZ/ZP8kLe0CDSGr2nu07Hh4u/ukyZXFd3mzsZdSjdhWt8RWs0c8hRNEgMGNhpBbvdEZsEz1gBBp
WK59aiq4aBUCfWkewtZCqGiWu3hyDLHMTg2P4Y/a9ifbnZpdCZkF/81yhJbUmHJipID354d0015t
MQ+C9Q7m5rhNdYTqzxH2pU/P8Gy1Ot8beH5bOk5/g1YrAiaDa6PmXcIMhg8XkWsh/YkOu/JgXc64
ZV7z38X3bwg56ZShdRJRB/X2TTLBy1BlnTYe4F7wD0saRtp7I1iNJwBIYuVXX0PXczZFZmbSxqVP
+IphLXDO49p0PTqDijk+pFUmdT4lVS9Oag6Mpbtj4qj6/TkuCAywe1O1jK327KXTSkiQ+IZ52Y6l
8tW+GQjTpMHDxBdasvl5xOvNYfr2QrqfaUckgbWgptnlDQYXP3pMhAgsp8S4FYTmpB3bwVon4G5L
XcLzhq5OhNp/0/WQ51FzTNXuPRizrm80uns+xAQDUJTNzGjrljTpvQE0TWICQ79pN2CZN+rTXKdy
zGznshh/aoarZyVhpCDIhBn5AwVIgHMKrJtRQgRf2i2G2kuAWdMTk4fz+qsmhu4O4WEr8E86I0A4
5Gm9RX4XAl7t5Ydn21kvuF9fjs+37aY0pUT6EzEGhlIV3LE79OVqqKYPtpfhPb34seZ8mkfkJ5vX
xrmNv4FdmbQ6Hbh6QVtX6bIhFjlEuAJTJu3oW5+RbajazCmkj81n9wmXvvLNzbO97gWeWieewicG
pqwzIe835VZrGmHFu2PHPanswx2AOhe1jH4XDCgAIE4KE/V30Zz1mcle0ZsuwkTiVaiBBmd3f376
joru0pUQBOUryUlzYcYA+AWPH6PXndxCule/U824plAcJQJSjaLSnGrrE5JuqY65W3WnTRqy3O9K
L55vAm5sRxZv+tSDJnAFlVFOClxjM8m4PPtFr364OFnLw+2pzxC7nwOTt33WIJTVhykvTa/t+aap
ZYoHhb13BtUesf5QoLkKbwWp29P1sbC3YoZLq9GK947poPGm5XhDB8RRH5dOMxQMSRreYQz3vu1N
Np8wYpRay/881EYL7N4Ee6es2VVkXcHmL2czJGn+Vwo6UDs2bg0X2B9oVXqFMZkBa41aermlq2VL
6L1/2GxzfnrFfb52awe3jDlx/NVt6/W43mh1P0CoDUJXkaK2D/JcWIBOkQVTfK/kzFqjgWcRKqvW
LR2YAxRDfqjv2STrAypKXAGWXdSPw4T6r/kSIPqemqL9mtUzzABIy7SOxgqB/0jvCabECANKGHGj
XR0T1KaUYYO4wf0nM6Odq2zb/+B+FXg3xIKGnzzwzHpX7pQDNzEm5zZavUhS6qMaCfNBIkgcRaCC
h4ddFJz+LX1vnp+BkpWAU5RHzx3LPEsmqJjbDFcPAB48JNBK2H5ViYo9WogOBZTzUYaYF2uM56X2
unv3pWCyjfvp4Beh2R/xiBRJ07gSqLmobir/2nNQT16vYv4Bt+mqn+7oBwwhDqePAeAIwyia5vxX
kMZmyh4Em//04T9Si9R3Ey9bjAKXlIRJ5VvZMR5PzwppQimG8Drj7NZowhtUWCEyqp852aZbeLQc
OuMDGRK6UbIbd3qMIz4PvJ6jKi9geO8dX552oY5MfSTafEvQ7/sV9aHAj/ZkEK3EHeMExSl+vzte
6Hk6aUUBAn1fpARrrbSDTOtK5zU4etxgbi5Q1KbBZcah6sljVSszoHQfV75Jt0UehRtHft3Wcegk
/CSiPGBuQJjDqDDVMjn7UIy/WVimfghvMuROmcnJUlQH/pxbkKzoR/iNkDgpoBZVlXkv42+ZsgyJ
dTATtPpLodQejWLHxDBjjJ2prCvrMS+4uBkkRVx5gVJEIivS27dzLqabYgkezstZg+/wB+jsMUFF
aS91tnpFXrh49cYXIh1uSp208oPRv4vOLcbsoijgxDL9LfPLo2xlqUPGUInB4r4Jg3zAMfqbA6RK
uqqD5rRsStL+mWpPc2uhMVxmRhMyuaxav7vccr0KOhtTA9uYZXa35v7ONgSsVUOvKSigiNOwr3cx
FQz89GW90/kWRAt+cBqWsmFe6vWHj5zJJm0jUAxfdzaHawLOpVolfwTX64Fk0384SI46YAsdXTXE
kmo6YG/TbGX050CQU+3tBxUoClWesKW2FlbgpJInhAaJ7pk9Bm3ah9ulCwmX/Lf8sV89i+Kd9jJE
1eQVSJUttlsK2qIVAmSSSuMnIW9rJk1b555NPPq22ZTGcRDovBQebkmnCI97GDzArMbm6psuQEyG
/8p8Tz4CaSxOsvB0U+tgPnjHMa1sLzy/zRJDt+uYTrnKi6fgBs/ruaIUeFIbleLg0ttt/y1oNs8F
pl8gbf6Nl9a9doZFhQIIghXhMFZDSiPjsRAbzaGI6saBMQQNmP4Efi9tCSdGxwpBQ3a5daCmrs6Q
frx5FTnI+xlCN6lKcyhu+Sc6LQHf2U+wx5FFJFK8fPT2P8Kl5AhIsiqC4bZYeKFY0oehlf9ahaZW
OU/R6/wvc6bXJ0Gr72nkjdNvFLiMjGhe7rve3fJJjbd19gaMTjyxeZpOGWCBoohzJnNtLHgQCSGh
jbIbT7uvVhDI3fNCLS/g0osRy67U6vDneWpBv5W9L6t5du4LxNBR7yFz4i0JqfHepQHK0lc6YI8P
rD1mLpoQlYa2QKBJKObTur2iGrWs6b2BsFG7NM8/vSX13oHutrHpndH1GKakdGmpJiU9GNyxMZJr
8aAGZzv0sUexUN0iiTptCD3/ZeGCd3iLoX+TVFmn2+U3K/Wb1/CFDCmQJ03uASfBClzutVYo5Iah
8h4cx4CG1AcHqyXqSoErPfZ4bm3arWloklvplT1xt0fdofZ6mg5D4CMIkmvx0OcIZElBYIuWGqkp
Q4XvnTLqG0luhVEH94kCwKbQ0sA1SzWUDgtdIxN6osOxJPRa5zdoCcPGUS1XwQf9Rk2luipwZ88j
lHjdW9CarObfbnOJrhKepMWy5xwopc/fBgfR6x8uRXmZiZl8Rg0qJcukUKd21119Dv2Dk3cbryBX
KJgdEnhjwRq+iSaNMmGVW/nNZSiVEEqzYELTFDo//+9b2nDM8hEXkTmbFoEjeNuwxOBJKs8cdPFj
grgYSchGzOMnVQyJs/z482KpA3Gnjrsvj7ca27IBUi0O2dNPQFo1yu9GgiUfC7mVLBuQlXuA+wss
ImHCv3wE7rcqHxp/7spCjqqiCnYa18xkUo0CqJ4FIVR5iotu+gU2UG29IQJ0uM+buR4r9u7EHCUq
KGo7usjcmrtbE4FHvL8cNTaM6AkmtPQQ6bsnCjEqjKPf7su1GmF1ZKHdVf04n0bM7PXMZbg5Up4J
0L1BXieChOWtrjZ0WMXquA890zF5LKbCaXRLXJNrYyXaZMhGYCnnpoqfckAfPDajUON4pshGxEiF
NzMg9IKgFLmELAC0DfubgJz3hgdnZYCYSuMYji+s/kbAuTEUTAdMFAl7dtKJGNpZWs+n5I13SyH/
+KBs8i3eaw1mJsPfhuDCcN7BPb30Nw2QK/NzaZeca/tjt0yoitV+xlkx7Mq8VJvmSgcNYimPMBzf
yze7he/jOppSiUykyBn/1r7DAozmRIZN5PcxmSiCEtmHUjoJ9FEhAl8QidPgfs1itHzS5FdGLIgm
5xsYUNwJal0KYIgp80B4xB7Ay3gbPlRczBHA+N8fyyuz4AdsWC0RRXB7T+Gf8xCGdcfWj9TzwXgp
rSNPC3G82nBS7d6Aa9BTHxWX7PurDUUfzPKv+l9Ny5tf8RSJ6s2AIFrUjPGrEyFW+eHPMqPR1zZM
BCyJcrn7CUWrueQEvxrLnhbUqmuQouLib56oYvCaXsF9RjEEHUAwM76e8EPU1anWSkCrMypiqyl/
Me+YwZIRBs6koKd4gl6VBIdWWMj+h9K6qZ26pUkmTBrBL1PKRTNeiPq9L57wC1IBKvjQ4uuOPUtq
sG0xsao6XtplCpWPjviDvuT0IvJTz5XDf9iOuR8ethiNHUe5dAoCmdEPNW7tPgwg+/Xs4ZFXR3RR
6KShjHTcjojgk6qPfEtWicjK56bu9atss5ssFThOrAREQWJmVVYPDtV0mTxL2yAQgd/Y/ICs9FX/
6/k/vDOBHlrCN1Q7Kp6jPMd5xcIIV2S09jQyzJ12whaPZ9ZWcrhKy6x5p8ykZV01+ahIArp7JkJC
+sVN8droabu4sOfYXgV1nl8c2zwTzKJxsRzvl7Xk98WmGLUSpKdryNZcYvSb2eFT6Je3BxQjYKvk
d4kgb6XgB6nqTNheSsmRyZg6oiHE3jBouirahABf5rUWxE47YMnETQETC286C1kXIfjorzVfurGT
sg5nSNrQuss0Y0FBG2ZQk1LDi4PePmxP9ubxFYSPEhze7XcmCtAtqz64pdFe+s0sSLhYyilWgQLo
hedaGu8FHWPL+0HrZa5d+0u7xsqXV+k/zV0dAARTFIy+q2KOxPkqRAPcMm8XgtqgZocZgONV7whm
x4z9MoU7OKqn5e4qdEHPqD46WFRocOn6qFjj4nWLsr/Daq6w9sAVGToGCLgbP3VKcn6t9v7NJE2l
PyImaJTPF29qjOM41pZx7hYryj+1YgdrddiDYCAYkZ/lt60eIRmrhbTzFj1agtkOg6CpPSt9DPXb
xpOzlwGHZR4Tw7Bpfpd87MjdBAyKAQz5gfSq/ReaNmA8hYB2DQx9P0bOPNscuMQpvebaCemInMp+
4J/tqRwA/DUabPihYeaLSQPj8RWM2yfnhpjSYXYvS565YZTxQN2ajJ4eXQKTQjWoAoNRWNN6U0Dp
IomAGzMEoxvuOdy1GVtn6Xf97Y4GyvB6RJd3yruYtFiUweaZl8743X8wiU50W/xKGQzwYPDtt+qW
aXHIsuee6PFq+SRpRFmmmT2Vt8t2byW1pg4U/v7Quz5PRWWofy2wjPogrj8B1FEJBRiXaBQqDAAT
shxCjRmo84e4woe3deqnIAKbWRaTT0Fr8qumfV46KiiBjdfJNSFDqIJCBixGRLRBPUos5cbEwtYW
1j1sGDA8ivKW9fmaeKE0mufNaEzVn3Bv7d8cyllko0xwW4jJCecL5f3Qc5T8dr/YRCQwwNLJsCTX
78F37rkyuVQeNgzYgE1jN/31qSmm9qYoNHPwpU/QmhKp3FsLA0rZg+uKw6pke8cdRJKgq3vmOdSh
aJC7F9BIodlroIis4DsK5OovKeeaKm9agPpjo+T5anrL21alhzQ299p/pGNCzASSN8eKOqneoRVz
93xUtAUw+pO28Yn9VhoMGUChIjLF6+ETMMcDw0hRxLnIgNm4VqXyvl3qrZ225bY0bT7M/WacwWoH
Wr5AON8opfj8aTMVV+jDVKEJJNMf+u9DOdYt73KjDxPycgRMdY9eIIMlWTJu4fK5MqP2PeojrfoJ
75QFlsS2ySyWQtR19ZYVOEXWMuesUE+Rvum4QFhbqvIzEFrNWxHNZlXcoz6H04x1fccPXIefSmyc
Aklw7dLJfH9/1+SNiQriLHk2mRCtXWBgBCQCMoYPQt5cloEx9p9+rRHAnBt78Ikl1vsmk8jwcPZ8
Xym130dsFgLautIw2/EjU0kSVaffxYCKbERfu84lFrlkMRs0YiRnCKVjRj++0FhZMyLwMnQnAp89
OMaZcQldVeF7N7eXBV8L3DWahMtXS/t3/EIB88iUdGFAZll4P5+w8BoLtPxRYN5u9FVqFGB54ZXP
InyriIRFm4lqZsKljZej3WeM954DPw315IIWW1NSTTgS+t2ixmjRYaHtE84NUgp2GtDv8McQD6ec
UDeZ71YxP0dzLgm6SqlwLwLFOzZYe2xBmD+o83wkqRuV0y3M00UH2uptUKtM7PjqPntcn7L6x0tl
gBQZCdB/PG+8vmtouefK2irqqznX0pqXHs6N6fDjrw8J2leiGwaJAwe2mT3XOcF1jn4DlLLjXWsu
ndEMta8Tur+66+JO7PUMPzzWR3vPrRWo//jqoLMvT9Vwp/zeTAHd5pUpPftS3bn1Ri+ni2nDcMyB
mOdNSznQmpRe5bfkvKHwddo+9pCJEkDHvO1mIudAYJA8UCK4AleC61Gv2YjFCsUR1mUKRCyV47Kz
DGGY/tPwxZUITuBlznBO+QVnF+SFe99U0kdScZW6bCT7LjKK8b27CQfEpamlNIpMZzymDUt4XNuJ
LhgHOBw4hnVXQIhFF68n789pW+KZgFBHKu9q4Fd05aWPN7hmexK9BvOvsvvdr7LHtF0RYqwppc6c
6HvnmZWl3GvISj/WrtywHwmH67cPmJ05/mREjbir19nhaw9hciSSm61oIJnSMwdgBKONDiOMZN0E
djS/ji/OVcnuXfLXyKnXdKS2Z3GQzyIWnoqNtqvgvTkWoRuJknXd5wCj/vFNl7hl8Bguld0NZub9
103yAMOEMGF2gUGmewuj14u/AuLMlnAIUB+NpltYkUnaVLanp0vRwnoEspZfM5HQ+bW1T0SJmzv2
7qBTxuHKjCphvBURldVOinIfU9ikgiEfaJyb1QO+Nioh6Vx3xashIg08XRWDW//p5pP54/zKZrrx
sbPzbcJPZcfmEyVRLDNtzfszEQIu8Hrnm4mFVtYH+XikLG8Q3P0VxbqZio3m5XrrxAsfFoV0+j+G
PgMgFnPpHT2Wib8wn/8TRPta9Fnk6Waj3eu/AnIW4yIF+hLO58njTVfIF7Q7ajvMqQaZKdI4GOk3
HOJ5X5pCNEv43xphOuKPq26tsuQm1UrCSDrsftGwx/O6yaFYRi44OBDiNfJYSNkDGVIcuyzl7Emz
gKn7nmQ7dpTTdVmOQgD0vcm7ODfYS4CRRtQGEGYPmJ+wZqsFlnCLw9gkfTEGMQ3O+7o1+3EC0Ggy
y2TfNhTqO4Cq+PniGgcc1N24AfWwy01a4NW3Tw4VMpPMQsILeGLfj/awPNc9z6Hr6wAZqq1WSZ+A
oSOxLFqkHLhHZOome0aijizZVbJef8tEj+1Jzv935/HYUqeyGnVYOZ+2w7bW0GHMcwHoHZFkdy2Q
FXQ8ZHxCeR3jFcaWZO+nv/++0eOIp2klEqod9Gj/V/UDNaN/2QkKLx96uNn1yNFHYEFLcA+HU19S
ui0xPjtXQXa+i8lADxa8bshb08BscvIINGdbqhPVYMMURPHSklj2W0rHvfhQvlGqYIuyxUixNytP
nHZd+hRigX/LDLMOy4TYpsJYYADbgQKU6wP9VXBxTlq5PsQWrlddC8pp7sJg2vj/1ungPs1/nA/f
uGkheaRWdiSu/DWfgFSsq5BS5odRz8qbVH8s6CFfqaVdv2VCPajasx+ayGNXj8xU6stsTTsPsE3p
Azdk1Op4ryIQp7vd2Cw76coGfXt4+4gJoMmHpbBpkhxnmZtI0+oTKOwbNX8A2LnI+2mAhX4iDGLU
5xoWdXTmoCa4GNMaEErX6xyGkXRSJnt0DK/tXm+8IG8Js5EU8H34P9kh47RhvlpcXgTDY92jfXtW
FOifqIblz0b9BX3LwcwXtl7jIN3Z+oeYsc5GFJ841DIXwp+MPFe++xXXqWR/ZGy3TajYD88dfl6x
ORrP7AnIV/GSlNiIvHI1MfRSx+6nnj/ounvkjMj/sfTb4OJuwqf3xRYfaJnDRakfyYXVrq8WTibr
6u/uam6umayZyvzJow7MpbdPsggKtGDwEqJ0P0KG6Y+tRVbz8FFbGcMcm2E+D201EFSZBNioOjeC
GW/34AbdkByAWziWLcSseY4NKdR1WiUHolP08seIYm85MKK5KRZr4TIAa3Jk/dh/0DhhV/LcoCZe
8v3NtiZrWQ0O5dce1qnWTUvCNlLVJE7aU7qaZfqK9jWg949/uMuI9blpnOW6MszoMiwUBlfIGkNe
1oUdEDjFCqQkefmf6dh1YzAexuJtqQ5glYtV8X2uafwLD1GFei2pW0o66FKCjMMOEtEr58fglY9d
o5IpsFz0TTQlQgeaaJSX8Sjm3/fFJ/5CTFZUa/ctckTqdvMU81kTA9FGENOCbQFZ/tCGPE7tEi0T
U+uw3SGuWgBymeO5U7bkdAN2CVVQZ6CJ35PZDuCJAwg6+3urg0xS8CSqUawA9yuFiWtJnWPibu9p
hp+xsE13OjN5OSSQyTiKF3v+d5S8Eep2N5egsUxZZsrr5MyYEMIpO4v9XJEcJSnZAmanINcQCGxJ
/TIhnGG5icgRsiEyRduifpUwJ8fshOTaUmoVwhWGNRGDcoEScLbYitah/QH9MYd3aeTMWe1UJ6hc
Rv/CCvI77U1//LGkcb1X34exjLYG7j/NkGfkwgbs20QhBL2pLdR7fVsDkIDurWjFqVPX6tr9fX29
4YS6DS7/lzlFNBkpEJjJ4c/czxpdoRnM0/W4JNjxtorFIza6HQkj9a82lh2A27oiKeB0/gN707jt
d54OyhvutBzEQK1f6H8qW0XJnxJ/dpIB3yKW17hX3A2O3C1A2NC/TzoeUfJ+e0FO+vVJK+ps05Am
YM7Zd84VCOY7gq+1nKxSZtys2uq/U75sTafVNDqB93ammzIpeO+yJy4j5nHZTBM+kYfcJliLx6Kv
J9MGBqaFvj+faAdzb03oIhgiNNykfhEHrfIxzYSUtProqfuzNQzUB5dBlYWBxN+lFdjx5SgSXul2
5Iyz3Cu4Its0UoTDFmJdakmit0urNElR9lF/S9OK336cvJuvmsZBvyaJ8LiMt3vvKbI7vuoQUEDA
MoZYvyzXIaCycDn9iRAMbZjrGHSDwsXMu32DWPYn2yi4X+7/ZKTy/g9qJXfjUqF/1SaaSoFKRCDe
ujB/MYazyZgy1WGz+ZjwX+24tGXquCtaHYf/coHI8/0H/MmCPeXjk+JbHNpESuMiBa92oaaz8MHf
3fqh6Gr8bs//S8a1ZfcEfS6x+OiAr6aVywxw5ZcKJx4CzCNGbKIYcK/WLelsYp5pUyF1x+G2Nqtq
27Pl0FHiQxmGIw24XOEWvd7XTUguVOR2MiyJU2OFXQGligg33Dtro4geRME0x2RryZmLHTdq+Hso
i9WLsmQFWauzU/4HaCUTPuzPLckNFWBma6FR3zVKghLV55LWudRaCct86bDuV17DgLPQcEySwkiy
j2SsF0kRcRqdzR5yBt/arM3bQP/9tmNlgFAsgEAUMAUPFhVB1dGEi/nHvQ95J6DP44ojmb5DnDSS
4HBYebNRrtw0yy0awWjjJPxEVOgdrHRHIKBAxdCIIkC76jK7NHqRQCV5BfrmztwpOYetpGMGGFRq
8mH0jyWRpmH5CskV/Bp8oP+nkVGwmI2pcFktNKBCWgu3bvKpXhUVVun4KqwSQ1UpgSqwedIf9rsV
fqOkbJvPN4hmSE4oVPpqVHMk8ubEhU73or+cX337srU3GFh+OQ35m0hPmTNqbIKI1DrGULONfisX
cx1f87vsAYkms8BbNSx/3GXgixXKapnt4wPJt0LSY4XVw51+B/McwSnhfRrA+B966zhosx1Lnal8
wZbfPDuItvi00Mpu6vZJ5n3+Z2REjjVg6ehoOXPcHzAVKC5fq3xGJm/b6/jZFwqu6DcM1NKUAHpr
Q/udH7LBEM+Nl3riAzTlxb829mY0jeH908MYyFhqQKi5Sn0o/B0xCZ8v7ASXXFo71EBdUE6LiUxF
q7vOhx6VWGgfYeIn4t/gmGL4MmFqvnaUQhe4JaW3dOcXjOIsgKQNWwW05+VrMsqxeQT15tNOgd2O
bUz52PWoXVhFv5pkEA33vkJ3ynHlBGmBrECkhALLmjMs9quPrwZ4rqdVTCoKGB0XxwxO/VnPLtac
d6neB5YKeINvMAUnDSS+j6T4YWQ1IinKpbUOZwMPRZyWgrUM4mduDbIakfxKsf9fNuTC/RX9GcOl
044EeUJ0NAB9fJ5tq1KF8dqelL3M/kHtcKt1gmtUH0J1uy0uTPYMZ0UV/C+TlQ9yqK4B07T+x1ip
pl1ooynlQwPDIRH8et2HTZ9a3QMjII1ysP+/tNkzRXK0aWUqVLpkkhVdMDw5mXWuqmIT1Vajv9Um
Z7dea9ZmUWlAAXBlo12MkmN6cvqcVB+deaZ7zBkknZ4aca1bnhj1bNFleXuQjOCwW2xxes+zBExK
7tGCksGMHePDyprMF0ZXmqEB1mpkIEIrpcQEsMb7byK/eyfSxPxJ1rE4N8Z3cYWKiUXvAYfZEOiF
1gZ7/8MlvosVIygf3TKoib/IqumcCy0OKmDH4v46rio4pQUN5wIv/rgxvtJ7/xmxCvvBr9SaWnUo
FhqnnyLWKcLv7+ML18krBsorlAWG6Wt1Klfwa/6blijCmko7Mk5iytlplDHEdEM8CW7PIpWw/fyq
sUgBbS7MyAle/mvhzIVBkrPYaapDSoEeQQfJWjJP75iZbhM5d2G4ueeMdP8i7/WRevm6Ogbv7c4y
XqswKLx/bxM6wX/hqjBcWoOrt+WAQbiySeqzrpgjUdheRphWYcYJOARGVF/PlB4oAZje6KF9Nkjv
1plXlZ3fd5qfq4rPFhvGyZGez4YK91raMP51Pc4uuWEDAQFDg6P/+HsYrdWyOz0xqpHzgeUE65/7
YVvXPDpwQbIOSeodGZHOJuYwBFREHGBYwp0NjUVd71XKF+MEwUXZ5uCDSrY/lo1Pi+JjBYjxMMt+
UfunLYgeF5rzivpaX8VHUo8zr1ypVs6Z7d3q6rZZigkG2WkZ4gBBU1kWKUKkEfLi1+4m2+4u7mMo
gFlco6iRNzeBMhVDnjSXvFbWV5h5hAqIY2cR0CMURfqbmDdQ2Vg0zGdna9G8dFz5zDRJdAJzdQZU
vCtjYgfwM4F3TU8HmwIKLQP+8DpRRQDl4kf367uKWIIv8jEginKdaEEi9yFTDEl5HKsWCTB18MQ2
gJOEzfUH/AqjpBJgl7HoiFB7goj675O/6dNiZq4ygWWiDrptocuV9yy+RXuS5J/97MY2ThqsDP2Z
0cO7RFev3v5DDqT7R9duFrOgqT2IoSok2quDxIaGFyuHLVOKihcEVZeLcEKx7Ug3EV4yL4ESj6xI
zIZjsbxqB3rJvKYTLy31IdpXdSRjwIyYfvhSDtB3RxShSRQtM28vmVAqFf4lkQAT8Adt3jQV3kab
H3f9Vwh34aL+c+FN1m8424KYArKEMTxqPYuP7vYcxgZ4yJ9jcLCNB2UQobM92zvjds39lGXOYTTM
zH91aUhBcAUjVyWN4laIJW9wWJd/+X6MSJO+6eQX4akCF50D7708EzQsZD3rdtWnsp0dZC4vdTtU
soEAvzTnkulBiDS1BRQejtUJ771pptHfA9AazRjh1scO8+gPyOA7d2r/seAGhV6eZt6lsto7sBn1
kCw6afpL58yK+8T84ZJzxRUCp2E6s+B0IJhBgZzhiydpcX9hyfTYEIQCV6+snm3cQGqNl/9ff22B
NNEuEtKtd01NXwOIHdqBUCuL0C31UkQIvQ1pd4ZL6mPfvHi+9rYvLpYeGq+enC0Uho0HI8ipgkbB
805z/m7brV1uyd0k6AWKF9xdCYmt3yudtxeu4BK58tZjDk5EHZcgswtRzVYNUyqcFonNo5bUUagc
xqEFUyou/hsRuBmmXaP2Zt/N5pUO1Zvp6F0rvrXm2Ny3ttHT4ttImq5th1cZ3lJta2wV1lKxlSAQ
6uUfU79dGItyTqbwSyePSCUvTED/qAldtfUw3kOrlsNQ8cIHhJHGJpGBP7LM5wSnwokfNmFDeGcY
AHBAQHcIH0g17ogPUtZlruo/VyUSnuxMDqEM9l8EnYuZmxY6yPFavjyM95vFNBDO4oYvSRhcRTbk
mf+SrHno74OJNu+Z9ti6AXCSSHDG3HKlyUKJxMZEZOPkAuvwHKMXSmG+C1FVgIB9DVDRM0lsiM4i
Py+aSO+s2h4r1f+KscTDZoslAM5Qb3+3WhmdgqiP0WBMPbtvTW6TCmhscf+JgNFd24xUFwyBaTHe
x6HxOtCDP73ZzwaLh0H6Hnd3d3hHsJYLLCzuQe8PtP4k95OXA4ZfKK51gU1QrReR3rXVjaetCk2S
J52xmWzCT/OsBTJFktPEGAmo8EatEWCSiGz9TGzVEOWwd7mq+PzPUjXJa1TrJFXF7AhPOQ/lbbpG
gePCw44y77WG3MdY6ugpdJnbVstv4M+xo2Ckbqb1kJ8OdaFpnqJY2vGE4k68eJC0OqIYgmOLjXgD
0CRwQvDvCFIxAqnWkd14jjGCdv0T0BGTkavkdUZD/ig3AbdBgvrP3AQaXfen1I13/xm/0aYSMunr
s/CkbmI5cICbokWus7wAY5FR0mQP7wXlBnjIjNtdNiJWIMtWPEJ+v/n/Ir40eLGoV271FqAmMX6S
B1d4cmOPY98haXDVvztzpqgCekeWuvPkTB56xsw89/8ap3B9pnjofRuSdlWMNwpIx/RuUS3Y8rYN
e3gKgs0qBu8YP9ZnP43Xjk29dAHEVdr9JMBVUNFA7bFAtnfUYsE0lBavwifT+hfpoMIxBjpipFKT
ZaUciBh+0lxshN5Tdk99s/c0mcFKDVuug4V4BA+s+cQKirGTVtX7JHhbIA7VBu/wYzOrCOD5Et1T
H5mVap/F7nyHVNIfWRVB4qCvR5e3COJvRKbOkegULTQB78/3LJgbp37WX4oHZqfXjra8QSP8MK+J
5GDpdBCKcBEOvES3PAlhXGUw6UdIzasipTHc1y/cLWn4dZbZgr1yBA5bSe5bYy/KcqnMRLKVprSc
j49dn59NAQEnW8/j+QV/DuOEqJnmCr+kL/1lqiAXUwwNtyZthl9cu28Mf/pX43FNvuZzH8uBkuw/
rnUuVuSB1SmfaktlqkHNMTOaMwDPfalrVb1lMMR/seyn01f1Vz6Av0z7uZDMeL2Jst3JQrBWOeQz
jKoHEhdqrOadHSDCfqa9AEd1yiSIQk7hC+KdSJqJuNpHVMN4z+/jLn490OrTQlhY7SlOlL5ajvGL
65RFAw8DDUSJpm375GHc4YOndHrGxeXhNUPKPH5q6Jdl4b/C01r/vnvEQMg5ONnXaYKGOZWWdwgR
vklFEcMAi5sawGiG0x6xrFK7KipK6ZwhiwErtY06TI0v6jjFmAA4ne/uP9QBMt2Wv8K+S9Elu/TP
24M7GHnEF1WgCu1XxSM89oN+SzkdTvoQT+OIwiQcJiP84bcRfBIyBW3y/ufhRpHw38O/2e8bOYRG
vr3Ldz9RAPG6K9i9KvMN9FzdZP1altbGJw+HwGwucid+jnxBBhIpudWl1D98PGK2BYg/cjAhSla2
6FT8JbXRL3CZ7hoHztcorJ769fY8DjFx2zDUShjBaPA7PuYik4k6AYY2ELZXcVT0Qo1ImLPkyqQl
kSxdxKKP/4DoInyRPbNAAed1ZrXSa74QecrqPbN1cB5FavibMg1ZKplNFvDt/Orkt6HFqLke48uu
sluQl504tsi3KVVuolQBAxiGFAzESlv9EMSFAiNlde87Ylc9A6jmaGC2HakZijb33gHNqaWRThhe
kUljCRctsRXz/ek5iW/ZBuXXigyM2tlk+a1XAMGEuAVdRI3m5p/ju8SVc5TmOLwO/U1nlhDBq+ZX
laaSO6ZVk32s1h5mFNoIulY1almEOG1v5jO9tGkVYKC7/fVtzUs5gBNnAyHOuvrVWU9upq/Z7Osg
49He1Q09I+3ryBFb98MCwELyLpBBYgKugExU06BT11Io0iT9f+nNNSxrQbRmBOY/s8n7Dc9cToJy
s+HbYhZ4UEpUfsBsG3cq3yws7j3Q6gQfK8sqcEFbNzKGQ2AbBo1QYgxTeJbMov8AWczF9Zx0//1O
y69tR9nsjbN9JB8rYmyFyY5Q+FZJj2tOED8kutCsrjOgOrGhukK3FAV8IEXPVWkv4mu907cab3Zu
LYDcLFELEbQZLm22p8H3kG1i+yRn7N926mgH1fJMdYfvdvBpz3+PV0NR69QTuODPK+mhCpgAUwP/
MFgH+BmikrJd97yUMPGd+YemDIhMvnoX+9D7ZL/+xprgvopYG4d3DvdWzr4FwGCBnvADclCYYWcu
mxIGvl16lAgJ0ub6g+OD5rLRvMpnq5P5CYLeYagznYpaPn/XzZzG5ZSeYM0xBzYeQ5FlR2V7fO3N
0bxyxKfYKwChBPfMDm9coMnsw+TYZQAvx6x6IZkp7WtwXls+2n43AAh/829qJQt43xw+JzulJuBq
mVKMZjCj7+Z7v+zGuQOOjFlvD4wNmg0xyLtPZWCBZ5Eo6rCjBen+ilZBwUwYEr2ps6xvIaGR7SIv
PmfEzAjLQeOSMH5lXB7vQKj/GBLxvXyqdpyD/zrLk/TK2s8v22plnOWTF7DLv5QAmYCKelM3y3qY
shzKbrUAiyyJ+X8bA4/kGnpLy4G/7YMUIFjjaHAj3G80uyDP9o6zY/cvyyMCp60dVUTEmBjHGCUv
8DxBCL1CV/cuCQTWkxYxJvnftAN4kI/fffxlr2U2PfXl+tvp1p3NOKAsFIizKcmYridTJrPR36qz
gtLdJYwePRBomURySlJB9ANReqRxSYvLOAQUT/boa8yva3brXdE4/EWF07cV0J0pKDEiiuvidb1Q
24KL55nto0uD+ZEdRV1YLLSLKng1fVQy4e0wCHiRdX4bhgu8Kk87ramiU46bdTy7Dabdzbg7uA+d
c7DvueuAsyQqFwBr5lVYysp4FM1don9boDq5Y0o5E8nvaqlOJWeSnxl/lcHNkIeHcCRrfpqGtqDB
FoJzBC8FW4mGLbtsmDuIv/frneHl8BUN+gzQVWQhOW7/uqWSg84uYXNUuqrAv9K94DQP7to7d7xm
ZBMy5Sk6NpQLYAFmEex5swznpf9JYzLm+z9yGpFWdlf0htTAXGGKfkyLO1EC/B2JnahmNYtxY/TY
ltzerYzGoo5oV6LL6OEd7o5QdWcI+YkZV8oe3YckmzfJ7agRC22H2No7bLBzmqKIn7LooT06rz44
Es9i1rnCQqgtkRV53Rc3pGrAstBdxKgkEe42P8/XeChFy3iElLJ8OTMKwipe5a6FtCyUTGW0LdR+
deP+Mk9JqtkIOiHUgylOivu/+Mrt3qKSkWKvPeGSYYP4TVZxioG3RcUbGHMddbhPA8HgyHAunHvB
CdAc63/Lw6FM1VZgQBU0UBu/yOxYTQtCO1IypnYqjPRaYhjlGxln/H2XjJx3mmwEPbCJXPoVxhX5
EncSIT1DoNcK/fh1D3w1rLoIspFF5RcAzhp0dL5cxXflI+jPmgF1ku05WCZ2NCtqZJxgaZWwhnFf
tB3zx+w4vYqX2i65WPY09TlRNeW4VCZtL0UCF/7jK+i3jTdVr6axY9K4lBTYrQbuHNQTJNXFmxpY
inNRpW8qy/mzN2GxKYEHC6Z7Otj2fysb2j33oMkxUQGbQMiCdco81LRgwwQ/w/uoRgwAyhm3Ytru
N/FZZNVE7ZOzm8/NW0kcKEAEXudx7vTbUi3ECvxlcuW47dysiBpdO+dw/BCOjH/cD/cOlj0efEDP
D1PMBGuyHxNl/ewQPSPZ5UtE+9F44iMkFu3k9weZ+KCUye93pffoBpSlvqFtCFFxEC/xxL0SOsbh
DIFdJ97DErzce8P6Z81fYuX84MzNxq57ongfiuJ8rGUxGQjxGDs0tPOKHa3iW39TqUjbFDj5qwmg
mmunLVVAT6ccl2zVPkrpr+DtBMbw3+pwsd0DncaqeOt9voljshztV2C78cz4NcYOwflk9iRHdWLo
40FiTJJ7bwwt4VtSaNAKWMctvVl0HtzfJb1JDQIOpDQdn3unbgMWufIaDfk5g/hTf1fifYkIxQvv
sISVxKQJUTKuhVxRhS854ubXQQWC7muEQEQNH2F/PwN3ZYSPKKpLTWQDGhbWLSjPVG6Ghm55B8sa
yFtmwWVa8Vj0WbgfD8Idprx58lC1PIubwQdwPUVOImAAAzLP5zI5CLbLlMNp9hy3ly2pES/Jx3oP
CC9RTWQNUnbfzQvyqDu4iEn8ahELg0fMqcMBUKMYIPJShAD00aGgbofFnyZDGrKu4/0cAIjBX7Wa
KG/VvgMIMUygxKDFp/u7dZOCErG6jyEVyFHLmKdb9mErVPTfgwdDZOKdPVF4PeacGB4Nr3EiHC/5
EREiLgCT1ar5V6c0uzfo4NeqquPtlOxUPW6RiyhA4OkzX9EiQ8WIRKtNV2NHc2v6QLHQhDk2idAs
FBL6QT2WljO6tLgVBVMIsSUAb1sleG30525/zn6jenR0e1ohPrVVUjibZOZAmFGyExfvJln9mb+F
qWI1iO2cXcJ8t3htPBcP73hwG8Dgs2a52cRXgYYjw0BYGm4DOQUZEOOHxkBC2PJqzZBQZUH/a2Wa
mZStI+wVU3VBYIvygPIcayJRH52OLxG726f4YUxtRqDuqPor5dEhB0/4N5liqQQ07a9YWHo7rJ7c
C4lRvRObthRT5x0wLN1wMwYRV8AP1TUNVCkzd5Rb2KOHnCzhIWkN8pI62C8eYSKxiy/k5oONgKK/
27B3DZGdGvzRvewpM7b+G+F6gnqDB5v2h4VU66S0Nd0b6StyOJlna/HyCF/RDLZ/UugImps/KaqT
gnA7d3MKWHp8uGzAeDE0NctubPThtmC4RrTnCcrWVx+hqzrntYeavxjMdY57Eend7j81Q7uPnVaB
iG0JlyfR6sJIoNzKczegNOA9wkxN4LY9BiAgFVjxj6N1JiQvkrSF7K9mumFraKt6mPme1wmPjRk/
Pcph16/of8SeH4ABZT/fXehKOuUmQbW7/C5OVX5eDrgRQjQJ8rCE1KJve813QUgJM/BO0aOLpAcA
ek7jNweGdsN3nQpwr0eFzrp5LgG+9yF4P2JXGGy70D351/PyZN9QA8DIfuqiMQsaiSkI9xHqZ72D
l80U9YyrlK2Qm+2VlJfe7JYQ/W0qIDb8v+vYmRJxG2N+pFv1sHYYGr124q0oEp9y1yCBnwaeHTmX
Ogc4Gie21Y1dDBBKqQPQYnF66Cr/sAeYBu2wWiXQPi/oQX0qwM4MzsfncWKzZGwt8sdZMWhKIrCl
j2dyP+xl7irS0o6//oPVFEhOSx2q5fTiG0EMaWea9LnTspBd3IAmwgxGOmcRmIOXLV2m2AcrrHlx
Mfwr0wW9+P7D08ISAjui3kJplIfekPMGf6tUsJbJAJd4S0cA2qedQ6rUhN9iUVfgJ38DBcwjsSd6
ksuZBfPZs798Ia3dZ9n3W5t3ulF+4SgPQ5+orbMqwLMLMcfJ9qf3cVwu02vFVT0A0cRowdm6yPnY
dzSx6A9vjyBLenbKB8vYHH4x6SBwFcsOdksvqzIoJc38ai47+QEUI/WcTL23ydnFXm2yD2Shc0FZ
UWJAFzW42y5DJPZHeFwO+hD5pV98ieK57OOjU7/juIy1vllDwwlyE2EKzjHWKsaCsCDecuDjjOOq
oksh7TrAPyABszRHm+DR36buvYtoo5xUTqwbEKZucXDIKnwrRnkRpJaa3IC3lA66iKJv44VNvPoS
XR2XuuUqax/6QW2RWw/+6dvizoTwS555MZrnaIeFpITPIGxm/pAVvnrkGKmcTfbJPtEyFneX6kc8
7o6HK4QI8VAZlY0vc8ar8wrpjvpjQS8hyGrCzzMs98oO6FANF2EZgp+I9V5I/Qlhp4b6e6bTPcyi
QFWsEo17a90avpPQPcBubVNztADe/G2z4BtkjcBZbl1TFfdfxxxyT4xLXyUJRJ7r3dDjdOxkqEGw
gqN18QyzO2qmVLdZN++WXB0EYPSAIDBxC8ZJ4+stNQNG3DjzXXJzltOmUCCEp5LkQCAzzrp76l/3
ufK64lSeIjHgLFHPmlA863xYrY+ZpHsm73ydAdOlNLEnZplP/l6/eSt9EDKo6d9GYFKXqzb6gUUm
rQf3FvL4hoThA1chBaA5eCzYl/imTeQ2gjjzU0RipaJyFI/hLLi1m3HJ3Cn4j1umgiGXsWTrNFam
3SH16LuLa/L4WdeIXbCNILZ+MvtncUM5uwFW9zFNbXGbCox1Oq9Ejtw8nLPoNxxGECpEzZEDQhsg
bBByPyXI6PaLDwYvnrB9ntKnrQ5k8u4gbFLsg5UwcjjjN4I3W/cMQBJS/HptDMhlQ1fPUqyWRK7b
V2dRcgdpzvzD+iUgYQ2t5+UCxcmT/r7/ntE68vxq5yDRXGmSLKLg55ShsAtS2FvUuyElXVNPjoE4
jVT367OvIPeGBmcEyQCOD80jo1QdVELdFQQcwVOG9fSL0IQo+H+M/nz+wYRujtYmH9Py3nFf5Bm5
7Jkyur1fTicdRjNHD/7pGfQQHalz4s9byrLpDoTvQFZti+M8ugfL5RQ1+n6EsJWQZQleb1vFwoYV
XGKLPYA6g8CsPJbamz05tc7w9yR498zGh/8KoAm/mNMWkFQvmI77GpxI0QVG5sICOuNsyw4vWRll
uDNM+5d1ES+hZWonwuzXLqIVjNXJeW+T1sodaK9UZLDhPQWv3eGnXtSIMSl4ZV+oA4SI7Spcjw/L
bcBQWn5hFyqUaM46otsAZQlxkm2Ri4wqjwg8xRFVvLJUzYZb+AiLdK7krSmZFYFMIIb95BpjgkyH
EWHAQWZjjgLgPEEgGaChL1F5ul7/ToNDeWAYLTwhy51qI7SA4FeyjOA4NYMZSNhAab7hwjh78O+8
do9YvpvW/atAt+7bwG6eOr6EDRotgDk4To2TmCJMYvMLmSVMFpjQOdzMmantzVqP6qGk8HcnMIwe
LUTRFQj9/mhA9c+Xdy+SLASZ6HhYB+biz2T/tR9DkVKUkzn95rh4S72TUSnI72STi8RfLWJ1Jn54
oUCWUL9I6w75ia9yPFsq7OS1IxSLwiy0UKgg3bOqonGFAoqQYksMr0NXreLSzm9WxN3oczRrxNcB
nGMm+rxenaZvCDYBTdrba2WrI2DDgMOO3+V7r+tFQT57bmFNB5W4iZA+PvXm46QFzQ2Ykt7kRrFR
cp5h/Z1FUTH9qCWQhBCjf7ZVbn4RHKPg16isyl7V48I433vOmyR1Wb6Ddm0C9TpisIJzIfzbWJbr
1ED62jm8eVqelOhKuc2B5oMldeOvr6jqRAYySGjQbkU6k1lz1KMKItMsz+7YhWH4lJkAFC7cJINf
IrGLiXf9ktTfNGwOv54LMC7KckNjjvv8eAijMfBcjgVMOmeJZdt0jdYQlIdN18IQh3oQEQUjk5K2
B/TVrqqTmpzqsA9kf1w/RgF56wYZRSk0tthSBC4saqv2b9NagxgVSeM5/mEYOTIQpgbtOD8cm5EO
eQELQWD3g/rDXArYfJONgLO/VTiYYX7wwXf5/O3bTFndTYJNb/YPq72m0bQWiqDAVbWdThSMckGP
q8jNwxuRIU7YAAzGU67DLQawBp5pHQazUla4+XWw3eZxp9gg5pn+ys/vZFtRlPqPYG1aZlJ1AVsw
aXSQ+6WPR+luBrm2z7RBbEPYq5F45lrKnRPyaYcgW+CXAiypx1ZkA8ubUllck5gjpVz52JaRw1FK
edl/onVnf5VdwvTjpLYVbaZ+YRy6PAN0ROE23KK3RuCKs/wDySYbhe4wMvFK1qC/EuAPH/RRyMlW
JOTW9ggF24GKmmd5+JQ3A6V2oU79KXljAKmBxAFzHa4GBpVAxbNVeA1VKN5fRTXQcmrFUSzXagwn
lcuuuPc2TSj9fhZknrznHNk3zoRWYeE7w1QaEVqA5AD+tSqSuLzSddvD4UoUJgdFXUKDXQxEm0Io
KP/Wrw7dfKt2ysmeIK1vRqOzaOiv0onu4vGkqEft68WR8JLFv+dPd3zHJT6RCIxIEa6+AiwjHlYB
b7gUGEgWDuno0QhyA7GWA7xC7Jt5WDRMTajL1vttgqNqY4nRhocpySPsu9dLfEKqLI0zYlO/4y8A
EG8ZyywGV29THsZb225BpU9kcTIPquI7yfGB3j+YZZxz5jP8JmHJS/8AJe11Xd0n9fmPExK0NJ6+
0tdnhm5TIIwId2uRTLzpgerK0mvpmoUf284XiO+hfOMKri6gg9Sz6U3CniwXzAwI4kwgtWgfhNuc
+K11bq89z7Yfb4vO3/+Twm+JVOnoeQzTe1/RMs25ZX1SshIDvZbrK+3si7W8Dp72s/uY4ujKiS9D
/pIyhyHsxVhsgs56EQA4PlP0+sFR2PBNXZ+HCZy1NGeuTsLDDU1XFedOdxisnuibv1KLyKMa90X4
P0pCVZwNzt6Nnrztf2oZ1+mkMZ70xt1SHCXaybyiIZCiHfnthkZvpVmPodYQ0oTQXmirnrR1hbii
htPIMHxAwe71R3QEC37VJgFs2fXPMGKyKSmfASH2M1pB/tpSrw5g+QGEsmdPQAY8C83b0hI95XuD
lE1GHrWds5+idVgP55HIlFAKXk7V2VzxAo86VYs0cQ4S+LVPv3DRpQMUJichOB47n9yUB3HQ1dVB
tNk4a4U//J2kk8U7BWUXbobQgYHtLH7EYMw46LBzB14Ee+V8v7OhoqKnteGmJAIZyIOUVgg93ucu
TWPyg90lGxiChwxkVNerhBcd/SvY8Ff8ctQE4IcxG3p2286NUuholmTvagci+ALsC0JDebi0TMI9
QtYZ5atOlNu7MgRnZCFjORjg12ldJOjxvTiqadxu3lpMf9aj4G1KfjxRYIDdS1v4sw4PBIGz0njt
G2iBJblJWtJrClBv311Cmwh4B3nJl88A4dYy2F0Isioy2sFqLwfnrc3fM6iIsJrcUMnIbmfHKzeB
CBuwn8LCN9evmUz4XrypHzJ54Tlewyu+GfLSBivaySk2vduQX0y0cQNCJLkgxzdW7xPglmHMHULL
L3c+waoEO9AiMvEGGsRSl3pNrBIpHNcPNcZZqdmyYkH3zVloTHL96iEC6Mt4SoTEtCnrhhG/fE9L
jbXyb1y7iLJd+M26laHsgrLpguZRZcYXQpf6CG7c7PRXk9F0EGrEqDj4gqPnE3ACznTpVauEZOCq
S+b4iM5M9aTecL+GJXJ70BpkvvfubrkkM/AlXeIAYAR6t0ytxk+i6I+41QWzzzEogEcIlAty/HC3
l8SwfDh2qWEkx4TCBlFCsBV63LquQjVs8l9IU5VW1aJ1H8bKpfVd5mnox8xCWQYbI6x/TUVHA3YF
1LlCpKmsNnG7re2jvTdk6BKwelpZCshf8Hxiaz8H/HYH3fxwp8PEqxyBY+MoTAWocz33j5iqa+dy
Fp++n6Pxc6p6uuLDLippTqVp/z7GpmfV8CSoU05SqsIAs8PhYmJl3vRuRgUzbxVMmO+SeizRlik9
5j+vUQKgTegXIcMmiPlcIMqcNniFoV1ShQH5DELd0OleOtISV5mQxDW9NBS+C66FUswnmKWC92u8
rrD6bFxoUr4oObiWPfN4n5IwRzel6QXti+o1jnkzGn5HrnGqd/4MkaCBtxtQfCZzzmbS8PWBO4/D
ofX9H+z5U1oBasUUMf1rforvUnKUlPvRCBrikdpjuD778D3LpajMs9TMgSMt+9rnbRBq/FhjUX0h
jDaTlxdsnKlbHgOvRUq/bjiKF4uH8uqCQkvIxPq8W0+YtRf3/q4EHmaFCPwrk0FtwhptQ5ifZwa+
yZ2ve9O9JUk7tElXXk4jPktIZPOvFYLZOp7xm+eN7XOZgIoGP9c7zMW5bbM6Pp24ko6L0M2g+CP5
GD/JRqdCUS87iEVwoUpmbzbUGXVXt5Ary8x9zlOh28TfR48An0Q1FxVGEXraTO2rimpt0K3KV1l+
z4jVSWQrMT1Mv3Beli9rKzig6PA23QMFlRru7LGxdnrr/DLR0/+G6/DJxYgff8fFdit54rFqfJT1
mF0Zd73w1bWaU9wHN/Lv9/OUuEygubX6poMD+ud+EnmQUB5JLEqr0PZnw+BXQ/UhtbR/hnviphMu
hrH7x3UuqvtEa/qhuqBWCGCa2LDR07Hr5jgPYmyrfLh/hPBBW/saJp9TAiYH+FoZOmzjkpnr6edv
Xn+lJ0Jsv/A7gB15I1YLs3KZ64vEhS02qCVOweUIXHgz8pYoZH2meCn9fFNFK6NOwhwC773GffS1
5hCjso2CAYbg9CO4pt71HOrzg8q6eYtZdJsSIS1NEyRTYhIzwdIDXzPscY6p46CLINUY5AobsrAT
EYICfvryoTlDZ5vc0rXut2IxeamkbDXbFICewgtbCwKhA4LXrwSr3sqrtpCrmcDmOZL3dtcgvnYJ
6rpTlFEZQUGkypfEFEQxCqJ2nAAmWXC1pzdoTIFWFqfqf2K87zmLolEKXMCjCS0ZtNoRZlmtNiCr
k0Fg4bLiLUcAJIY9O6mmlRsafCY7cadWp+T1C2zQsLOiI68UtLpAPZmftermstLgE2XPqpxL6bYU
hPkXcTlAZl0/8ruxzLRNTAoeBDQLBntp27ooBoj9SSMKV9wAoV/HsL8utyQHrJpGsURCDOT+VabU
1PWg5NCg0XGSb1/Sc1Tfd3YdkZKS/pt9IsX7ylBCOYJFXlu6Qb4r4DYxNl32GNdmC8OtDJUsMNqT
wKGe6CfX2mepEwfJn1OhHoK0Ig7s4n9nJ1H5N1+ZFGKtRTRPdX24jGm8+TlbHQoT25yqOXIgeSC7
psIvNE37Rg4GlNAKJv/U/yfzlkOUjnaobifYgvJdZMb92n5fO1lxWDS3wziqCy7t7QI7zGC7BykQ
bbgc5yi06/jbR2hfzFzmN/nc1vMVBHapFkaR+ptOby0fLMxt9LGgZUcDbF4YhgYKPLm5Jjm8VlC0
OUlpv1pNuFggWEFSSlSn1zsaFbPRi3HGyg3qZKy4yuXr2YKGcd+WfYtLyXk7UzS5yktK37YcnwxF
48XqVDOoxykE5Gb8fIJB650cNYv0N0yEHF8SeZLLJoKxVKHzD6YlPgzbBzpf2DQ/6mYNQPSfmvwB
i9W+CkiLMnBAzFj+MmsOwLvnnOqhllDG5om6nBW1LCENmFLiITFJCFHtg0Ga+ZbiaeloJwOfuykd
psz6LTgo395RBFoZbCQTBQV5XYCz0wGfbP41/T10kilTVxArep4+n6OgVQTtrganLIBtyg+qsxsg
Onv244CJrPZR9CsfIA8vZpCbOyOt29rcrQMSxKHz4tY4ivZyu2xOXkfs4YSodJ2DPce5mVmkhWLp
zQx+enmeuKo0yzbYBfyUCNnxrK0cxWESupQ+GeOS43VBTH5sGSvIOEvH/xccKzNC6usnYAZ9c1O0
1cabYrHEWVZcTre8l56KnrUqoOnlvq9eQSIcWusiqDzRC0ad1i/TcMUwHkgzYyK57789ykrpFbEx
27zBb5QXykmO+S+PtEvbUuJAhkRodSQqyBbviTlenkbJWAvSvo1JchFvngy8x6Ojr036kGFx4GOV
VGiuqMfJWYtfpn9JWRthwsjNlvnb7NBh9bMIetOtJV6xCRWLs0wtCtd4iN+4ZbXbkkWqh7P7PaSr
srQr12ayMk/bhuylIy1sVefsDfuScViZvhHgX8i0b+OrEWw5SR2+4C1Svjea0BvNgKQ/zbSGokKI
bxaxXtsLIOqD+GrAHqg7iqo4ydW8GF1oIH5OJ5Wao+/V8huEqYejJP0I5XfPZENxLKN1wSmnHBSg
DBtMXyh5mg4tH5Va8tZRzyJZY2EG80CAZx2uMp80VAlS76ikLkaf3la0O5lB3tYL5lttbvON1DnI
41U1MW6CNerwEybrFQ1pXa0j4b8Rw0x1azOpYsCIQRuQiJD85bwddpxfaBhAlidCn8ZA44yk6Trr
BcedsJYj6oa4I4WVTVDGCY0Ix3ekITQTlZOudr1daRkXDJXEAXOVWA7UcTh7HGnjMSqcXhSkyXe8
cVz9gr28h3cX1/kmzPUeP6HZiOkjgOrF2A7SeJGGRiRBb9MugWpO/3VkvzLGa1s+5HhoSMsY1aqV
ry0N44nadTwJ0sFGhvAhvOV490sr8lUpvvtjip7/VyvD57tZ1r8Er2u5CY/8lQPpAlPs4DN294iw
dA75axUnwo3UtV34M4ddUoKjgYJ/1Ohpk9DXBfdGKHjgddmwgaa9fcunVtAokLRq/kkqxyto5N1v
fl0YIEF33Cl958+uMBfWb5huoHZ77tZXNovvIZyudHh7HESxdahaQZqtMKW+Pk4MTRiQXnU0UGZb
E4PwCmRRUS7ZsUtS2mMVMUfhRo10LlR11I7GJz156QZBnlQD+PIJajKLwanHCinuy4wSup5v67yv
jRAzcR27QLbhnR1e1UzBUw5lYe96H/rJcAkgbTQcK+2IUzGINgzawmAm+P5RPwK+z4C+FjZLMz7B
gsd4BZkJstOKR3c6CqCcK8fbvaRcH1xCjF6DO9cY9J/iHc8eadjUfke2l3iadhvUGI08M1t7T2JL
KxLbxFxSZJhI9++S/5b4zasdF7EyrW1nmFjVqSu68UIgt58xfj1yUQ+3rJ3H5vSTSqnZVu6T3znO
4fM8o3dWKk5PXwr4sJAnfm16k8nCmEw2aiM3w3FUZf4IrFf4jtRn6zpEA/4XcNoo5Sw+XwKJeqeY
9R58datJDLR8Ee7AIrQTG5K/Vy/X6qWDEME6XdKgCemJtKr47taTFwjfJEVg3tv5Vmn03aIoTtSO
6wzNTC6vrRl7btv4Q8XqOascTQNEuXE+mLW9EcYFr4NAh1D4I9+yjdPcoIhPn0+pNHjSVMHJuh1F
9OsdzPNUy6sE5yGo+0fJGSmYUaT2Nof+soiCZypaXXe0LPykpWWPcIW4c7mTYLxW9fGSUjCKO0kR
74taysCbbNR1uKFZTa4TMyT/pDcZEmS4HKORwDIZXtl6LYnWZR0SppmBivfDtWM1sy36Ub61AZVH
3XDX9UXwUnndIyxyDSTvN9t2Ezu7RaPRfFl4+HVQRLAOcfePQ3DCee2djT1vHLylzggsHAcpRbdX
uw2soNry7zJR6OndHUoVkcWqF9XywkjhQfH641cGzscEKX/8wQ1GqDltjVOVEa4D/fHTkOlEd/SM
KPvuqjHHV6X/AhPlYqLZoVVJUhzAeBD/IOCYRXNCgMeODig4OkvFjsB+s6kPt3eob2YiLVYZxv48
TKhJtCrKJnMQ/vbXZu9kbjhQdC25CVhm0J1o4CIIOQl7M5f+eO8A66fb64tXo8oaFLx/oRrwuUDJ
W5DTUTTrtU3suUIhd4frTbwHyNIKyd1krLTxWI8O5g1stIgkHl+NI9Wt9C6DF6DPzrief2ybsmyf
MYnw+/FZZqADEVIqeLSWGQmDQu/+jWDL/xXuQEFFzLjZvekNXse0+TGkX8zNsjSTGNVYngztou18
0z47mV5aP54QAU4krY8ngc9FXI6UeB/546Xpj9wlB4YodAQ6MJevwH2zHGPBP3T0KtLhyktVsxhp
mtNBD+V/WUkanrDewfMuTZNGdCP1iVFZWsS8nPjJ8Q5JZ8D8T9MXZC8c4nWwXrEB5rt2HOuCAyk0
tjaFUBXgNOZ1GPX1mSBqPtTFN0Z4gr6G5+ZuwROccCSwJPNrMyetigKm0/PlDuvX6fgqLxuonRxm
AnhbRqcgVFgUSd+RMkh+WQUnTD5T8HW+Ek6FOjy497koHU4YncFvDuOgoZv7sW+DFsmH6kVFqQ58
HsSGi1tYumkhAOCPOvoxyWZEQ6Ls/Nrny9CzL1W9Vr+wEbB2BQG7MBKuPRhInL8zLTGNg+vUEo7t
EpYfJ+M7IRQwh8HVb6gOuylK1UuNM38es+nYi8hUzJo9q1mZfbIQNyULWYZNPDvkAP2ZYPZYz8OO
0o1sSldauWlltXTqBD9KWIDEmYGP8qBVX61FmM6TKgG2KG7ahR2GEOqUQPozGajRHxvAbn0GqtM2
bkfufFi91lbrVp7u2G8kkUeQvUJkc7wnW34xsUGNbjYVrbj+is86xjRTlEBZhfD4haCBmihXFHg1
KnvrtYdGgXpW+/TiV/rpZU1WAkwcu95AuuFt+bg6SxhklEIOyZRaqBzN+LIe5MGhlytwco63h7ty
1JQzgeOKGaAon22wK0fTdMcOk6wwFKOtVvOyePMRyRVi1sPZZUnay4SxJDfXz2AR6xX9XqkBPbvx
m1vAQeQrv3XblrOTea1/XHNQtiUxbMn9oGEvYHd/ACbysmBS5lSn/c9+7FnStfv+q2H24j7uRLoA
mcRsETti0C5IZ2dH86+E3moRpRIlryzX9c1MF+e943xSej9xodpWJaf5qxSTX+rs5vJVtYtU3hny
k65wXpfUZ+jRIdcnpKAm4F6xW6Vifc7lgfOMQQgJ5KpPEzqEztiaLsoxJqvBgB542xOBXYufLid6
F5/FQ/KgQNG39hUxKr0Z2eqi0HVwJgeDHNYq3+aaeSgO1/fARkd25ArurU52uJ6rTEP83FLIQRWn
ByE5W4SuAtI7cG6JeMKUmT1RzpbFysFfIhDrhpASgikwgbXP+u+Iuct31rrx0UK1QiJVterAsh41
QG+er/PW2fu+qSgyB6WGliTcaODImoKcPQfKHHr5bwEfgzmojWAeKbVduy5zWZcv0qqnt/JTJIhO
OfZegu8YqOXbrBrbDG4WLEEjfgTkOO87LKxdA9+GIt78eKP1mswadA/U+uhgDvcazPhUdotATCah
qJ3lhk7N7Up3/bArGzvIk4igQmr8oG+ZnXL7KbR5Wt6hPWGt1osrhlr7sxQN8j4uLgC8JCdddofu
5ZeSjj7tgmwSksHi1sOlb3RlzArMwQPLUcNJ4hezsAwheqMIHwMtiPp6PFTz2Hh8rZHfMZ/MNTej
NbUw/vALiR7jwJb7239sXqsfg+zrS0IOXbr5Lh7PG0UKB2BaeaA2cXD0WMBqzeOSQzOGds24XYrN
bpQmCrMXkLxWPy5wpLcoqjRQ5QkC9pwSouEAS31SOhWIbZZWLotn8m8i154rt7YN4QyUSVfXieCR
Z1XzET0ssBh2cD8n0D2vaqEdmbSlfXX9wJ66JNgv5PFVlUAr3OWpfTz/HYrKUp5dmqBdbUtDxkBM
e4IaJGEx7f0Nw+EJY8O/P204NNSuiQOYxO/kW0UrP6gdyQ3DJ51b+HmmtdEoVqa5UvLQCNqIiBnr
IgvGcg5sV014t3oHBOl3eDXLI8+aHx07s2BA7zB/PTnQSDVNY9JMPPF9oNeBvpEJUw+w3Qsr3H8r
GoUAicCWAinQ5lB8RNQZa+AdNmVww2HeK/DQGkzQ239rJteCiaIHJdUdzVKM6ThtrAILVUsWfJ+S
EBHeoo9ZDL31d0b+hyA6IFvZk+FcHRNXF7E3l2WuUVzgctcdMJimmDb1s9YH99zeiK8H3R/08WQ2
TUonZ4MpxZcFhXUmlRxXKAqR/e3QB2o9nuEF+GUSrFcl8ZOxvy9NNpiO8z01mfjS+bDPgqXLascJ
zGVMHaNtW3Olc9uCUXj2i+AJCSbz3O0ZDSh84UzWcxucumnY8x0Jo3+zFVUNMmNHB7WD4d+CdTRk
N+w1Ea07qXmmews9qvNrRxKoz72lYlP6aaahKNVMtAqt6vZGvIaMe5Xp2U47FrjO0l9wdWEdr50t
Ads9gYUCUhtV/j+OfVA3AGi5JDUxZFY+iuFuMK5XaIp6za/pIF0IlJfGkkqPkP9bvvjDobuQlF15
YUh71ipnREDI5vN4lT5xwN/VQOLpP+LEMOdtJEQ0orB6MtMQGZb3lEBAmUUnkOLYEPfxvAVIV1i/
d6fk9+lqLgRjGEo4R+LYhq2A3A2i3PQGRCXw0l1WOXQqtRCxUYOVswMbjXYkJiORfOcmPVS7wqkn
Q+TONkHtGBUvyJQ5OngpBaMc0nx1Ytf2RN70S1fXQb9bvfx7zqhanGOsnnEU4TQ4TWE9MI9bgwKQ
0OD11eS0zAjYDiJd2nvnnT0W95hABoDZm8/YyuIL+qpLWK1pFskRUc0dplPuMD6IPZ7EB8zBUowL
Fj9uIusLzSYJLoXBQtk1mi6sAhBZw3a4Zc0Jtktbbb/Vhe3ArTrQPEAWUwai0NKj4ZiN4+cmRZlF
37151Ml4eNQPKl2K7GcbZLSmOHoaJA8GQBDFx00jeTqFE78861QyecmY3wxrQlzHf1OcMJWZhSsU
UIM3k4+zIWOOsXnzpwo0ZfIJCqqwF/7ZPpR2MfJwZif5L8cPPS5R32b0lrkHGjTxNr8WyswFSdyg
OvETaatfKFyaR6qqQiolFMnSXqLKRA/4bWEOMI4zBftD9ft2I5vrioKEi9Y0gsbHzGJrU+dprVxg
HKxvPucZfNCpouRJjp3i50ndQcDtqkd6uhxk/QYA02LEID2y9Y3xJ2Q+ocAWEifskCZJDXv3HU5j
vOJycp6z1pF7gslqZge1H4cnQHbFEuEI2LtkILRAUB8sAUpzkd5m92dvrUkLFWZr40w7xv0zKjBx
4U34j0oSXWYqBseobuDiXmVz1QV9hExw6OYvNC64SrJYpdsWoRqM9TUwGE6UlFNhSO5WwHk71iPx
8QMxKWqt4iNA45k4WLESCZysRdLu4WxIEOML7JXFdH8dMZRWoyu2YGzpO0TNOkjS+6xMvAlBeLNX
Le9WTeRnRer4d2eRJOvLSzpVWfTX80EDzRv+ndyyfo/VxoQ2Jwe2Guy9Y1aAJtg/hztMMA/bFfg1
zTQq+dbpD8k6TT/gayLluAixPUdy6Yyec7VIAnC45BnR5iAIsiLRXfx5UvJOtPvkyEWoRCi4zBMW
TlPExKPEm7krRhLM5EqVrg8nGG7aDHQdHsJ7UtVBOSTOHD5vCunmw0EAKokx3bWCNKx/4M3lERRx
mDGL8KCkV/jSmsB61f5iSW4f0phobATIiQpms1lNbbxGhu/3kANQ/gs+xvwfskgPA+keE3eSLlJl
9wFABfIfEv2BuF6Krg8w51OiSdS2Arm18lwwG73qkUc6ZfpQnxLdbFan0yOsu1aroW6Cv3CdgBQ2
V2yCeTHeWWuRf5eTAXjrb/43I+s1q2//uDN1yMLM8ndy30XDK5nzf0bk7ftr/Y8+z0UdlC1cAqjt
8ZCib9G/hxhwB+2ZbmXyT10Tj+wi93RRRt2wGcbwAQLpcEYGqTIvEVdnXzY8a2ILANItKMhtEpr3
e5NDOlU6thw3OLmh4WaYPeTCkxmGGLpYQB9ePy4TKyZ99NwYWN4wVsf1bCK3a9NHA3+5DEkCJB7Z
GWK9ub62JErsqqfEn5IFX34td3UA0/1lO7h8qmoRKl6P9b0p9xfaZH0lgo/tYxB85+r3OqMfCUb5
/HvRsK+BZL5F4JPXUbDzy7LVB5BdBG82pRPmGpFF6eAHdz3fpdqEDIAkPe8BeNXLCDIe9x+4ZeMp
3Kts3lfsUtrqImJ58PXEcZvhxLOW55ejhn2mn4eu/FGEPVYchIDAOKYoUAnl4dI6CE581ojsmxTS
HmJhINDNtfsC96r2v7+VQG7zt8X3a0NqCPC7tCAkPQeyMkuojC5e3AkAZI4U6sMNci1zZtaMuO9o
eSLgo/ySoy6WCv+2Nth12IbtItRuv+hNQJ+ocs2o0R93ZWBaVpBv/HS5I/zcZX1EBPMwy3LxU8cF
Ko2MSqx452sSPKvpLC7CbyclB+Jn1ORlUIag+YFTlErA9Nfu4AmelXMApbUfNYfRjVog4YK8Lrzi
EKCzBE/1wWEyb5fDuAWWesi3L89sZRKX7F53wguiffHcJ0Wf9AG4N0xAd7t9pU3tZYSgD0bWL3eU
9V/qdX76EogrdRAMZmMbsiM2y3+l9J33Lt+yLSFBUjNuLsVMnBAvUPXuTTKrxs80mibQUUslCYuM
0GBALTv0XBTW81emQ/hPf3Dvr8x/ssXfhNRDLhYavrXz/ojGKcOVY8IxMCvaCi78LqdN3AlGJ0Pe
toUcNtwHTg7nLJQ+un632i8QOZPmkGGNQOhJhzR6ujhdAA2VpCRDrIU8vDJ+Np2sAFRVwz3fXdcf
4akzfcJeYlOKr2xZJNXznMkjHKLkqQ0o7oQEF5Iy3ZCFp05rZjXp9IylI9dfaCFWPXRg7Tzkgn20
xV8iTvqKeRzoqY37oYqt3CrjVONgwnVnhH8O6daw49EFP2Tvg+M+DtVinmCUZ0WzX8zUCB0JqiGQ
DD7PZqgJafTYeP4fiVbRP3jIqLn+lSgxQRid2qsZSSh4FNmzF5gfalYoN6kVPcKRFC3NNK4BVZ4f
tJ8D5VjxjWRarz28zfXXvoNYw/jMwB67TH2MveEWSFKGod/MJQn+4+cE0noidoReXmAFzMUCINBs
0dDV5QU7jybsBKDsi7tNzmCLe/ejjR5QTzW4uB3p+wPS4qz5Pqo1360Ervz9qaehFtK35VZ1hqgS
YuZ34oSHVokAjuA4AMqCmFoWTyX4xfkCPsUaiBv6V76ihPSCRw4w6IPVsZ7POOhXPjbdEkx76GVb
B3EIJftx2CbQBbJwO0+7ypW3nNzfzc6nrMdDyEdrwkowcGaqUH7v06XvT+svjQHN4AuNdcRD+yHZ
QjFKwWm6kcyR0o7QnDg56jzfwGF+cNmogOrT0pciE2VGqekzSMOjuS7rmB/SHgS7qFm2++m50Q1e
rSRp8tcdKwcJ/p/RoXsmWrkRl9YtL8NuIt1K/jRRZImTHq6VX+O1ZpptFM948PN7mkdQqTcej2Rf
ZA4MgnXg67KYqVp4vBwbjbSFa+A7iaIv8A3G6dlzOU/TYNkqkrAR7rcsan76/bL1Lwnyj7TY6hZd
bQ+sD+nIEx8MSmVL7Av9cbYjRp6ZU1lbEdd6utk4BeTW4FfOQSSTbLz61hAu8b18BJO4HA0abXNd
XaYOnYySCJLs7tfxF00v1NLGjJY+Nh0SKMsasnCLMRkfaJyaNCZaH7/qfEsPJMzLeEWorbWbPIO3
lw2dNYToS7uLoOq3T8cHNIX1QxW7Xv5byy24VkirfOKAX7ZdZjv7k4gVJGGHg6tH57CiZ8wyu4y+
yh4Eh5nWnzDsK1BgPG6T0OXq+Q0t+QBg6DCRJEU3cu3QZ7W6ayg2Mf1eySUWtlpJcXx8hvsHaH61
j5NMBHAUdeIN26w2b7VP8i7V3wtxSIpZVlpteQF5TAhhkH23UwR3AycpOlCRXA6aI9XkzEiSd/nL
5bdoE6q5480rObHBWKptbXVlTYOz6NSmxC6b5j1ZCRU4hx9+oIKuQbNu0ELh9G+XdipFGV3wetBV
taWXsG53nAAZmUgcTCz7v3NYzQ0oi+o9K53Yxr6W8AJz5xSPGj5QGjI5YUxPJREp01oqhCGHaN99
/FaNVG1HITv6QfZMpYda33jSd7u9odY1pPUIThL5ddl0I8u1BFZygtwY48FEBo5YX6K3eXHqDziY
uIs6ynwRgkNo/pFXnL28TIvn3aFYfjyPaicniHEAdw5VHCv+yGjbv0K9zS/bWl9ILmIaleS0D4p6
MqVciyIKlNSHap7lg/ObQmSv6QetkK16zW9UWHQY7C+/zIj2mhtsyJtdquPDLN7I7UKEoT+e7Ev4
8N6RJXO0WWedEcxMzGZoNP2TWpgj7uGooRjpjDHU6YobAkfszvnfEptlyHwO5PpNRdEkCABj5CNS
4gCQR1lpHFC95LK5zwn6E7DYq28NIMtT0ua3pw4rCRIgFR0rdaDBIfGbxQtrxfvjTzHHcYgz3uzA
UYvIsMgsYv9NO/dNGQ7LElmf4gzE7eWZ9XsO03pC7XZH4cil1SDvIjpfjRzlSuigU3/cauTUhWBl
p/MHkjPOYugY5OKoXLzrDGD5//CbpFrY2WbzmmJtpLPpqMXnUsTYJA75I0KZ6ji0ijUGeju7qkU3
3XhL+9T7L50XN+GP59zaNJWmEqC+HM0TLXSvsFwCJC1MhXUyZQdtDHjfXjayN0zmfAW/0U3H46mm
SZ8i+3SDYHwBJgdz9HAbPs8667zpLjmkMJvip+twbN6Mm6LEoDFE21j5m0B6+NCcst/rnw4ha2+Z
OfgM/7LQPWiA8EsZkqxVVbIaQHF6Anv1KTGvG4gxCwgKkYyTU9HMrN9aXfHZvXHEqMcyx5kyCkrL
aYhASLkjyqOUMMafdldaK6Q2xUL8D+xJ4VqLpCH8Ks3egkO3vRZgddRHJSxJToi/yk17UDuOvYBh
N+OcpKyhWqByjQwGdS1u7FfjUK7FjM6PuKsSd5v1BU5OnyHTQGfJoXlIjMEM3WuXdjBxkQfNWatR
5T0TcBNYXhUWpvxuDfLQg+SO+JdPTDd2hHu8i+O+8P2KyoaS5EJ63QNUXNgQ1tK/43lTWM5Y+h2D
TXwUbxgSvweyCqfM+R84ReoW9Scw5GKZZk/ju5f9fYIs5l7M+kvOIQNaLLETX2VwJ96n3FRzP7VY
iH6h/jZ5EUfZRZ2nXjslP5L2PIxf9jjPsMp65oLq2fo8qGtGJAATlXrwmBLjAgdOOIpObhCnwfT1
Pu27OEMqGsH7ec8eFKPEM2+gr95erBZllCCPdxLU412+Y2ZLlOv3HiPVZw89t4Lv31h0cYyUhkSn
M06T5Jw4wRsm5npF1kY98JG9ZH6HlTBJOn33DrA3VZ9TUQ5mvB8PkTs9D6n1JPiWt+lnbN5NnDbI
7Xgym5O1qHRJexyCAXgAlkI3mfIQ9crw4tgf+2ri2PcALmxNnmL/d5ilFrMsCf3h404BSUyK8hE2
wOI/QjsYE+TBjEu6g7Wsrp/J7GfvyF78nC0SW0Qn05ULErhPMvAoi91/fE+inHOZnoA16U+rqR6s
+1YJ4zR8zWNf4XH7EFH0zqeiSqa0gEFevujA1KQyikR5yIq5oC/+bzNjCp9Dp9CfrLufCVcYx9B3
ULllOaXfxCKvjHKWDg/UxZ3I1CJBOf8le565jCW9VT7NkyqX7eHfW6n2/HWaBlzjlSXJldXT5Ru5
OmlYgk4vMUEHpHveLUS3vWfzk1pEe/2PMkbuiH0WAichwhV3l/Jg/5ENfl+3/g8jX70Yd7CJ98Zp
saYnZks7Q4BVQ53CmLTZjCWDgRYkRhGaCsaP72qX02m83Q9apza4VWbfSyE36vHXQ8YRyoylj1mD
4xqydtou1UcD2dC3RfpePxH3IbzvLq/lwQNfgOrMGOOtaUJJRTQC9nXzLPtev4fWB09+A+ZmLoyw
gj7jAsBBbB8A/G3SaxTdGC0hMzijSSSX/1mANW/K83LmWRXsMTt1YX9EQxxGpUAKsJpgdub1pdSP
JnNwel6lhm+OVXWow/DRdiFRmufiw8xo6YIskC54zv3c5HI9UQwjWbRWbzbDveM96jn2XQGIvtK7
ghS6SvYUMo6CkkWerLLlrhOATknG58yDY6vPU7SV63H9UCugkVsJcIJK5RWOKUuPPfDp8fb8TGAe
2D4yiLxwTMgQZs/ltpmbTeQuF1qyrfxRAsCEW4Xxxw4NKZUWas6OvdKHbQ/YyMohoR3jDLF2qrV7
ieQ6YVLU/O7SBC/b925kyOGBIH6XTn9R+7JnG2X+qIBH7k5KYkpSV5U9HJeb/9xBgYyMtpkogUit
SD0t5cVaCZYAEfxSAoXLyBBBAzCdRMM3sE+3Q03CdOvAaGh+um972AysM/PCFEJXUTwN3spUkNjQ
BBHv92kTDcrF1n1yCzRxaUNclACPNGZte6mn2/Ws4xZBFYpPbcibIwYQlqpUQQyf34GZp1dLfeyR
9AAde4vVJ1pC0KTQ/qf9qKqN1mXGGvlOOQuxeHZ+NyIpiAXtEm+6yTrw/Lvt8aHcEs+Rn/h4FLbk
RFrJDV91Fo8+yBpAfmD4CObVQdd0n1H+VenBXsOeGrm3D5YySa8dD+FWO0dseocqPwunsRT1BcTk
WVa+MwYpAXzTsas9cvWpEXhKNQZhmzPtODMieRGzYVSfGD6SlYrugfI2ENxK+4/ZgSWMiw/0BN11
W1EoPebT729BlPXdqPhf+dmdZSXk9a8xdy6IXqPQ7st3DMuKitEeMhBA/j8EVIFiF2WLhZT3fHOU
qoR/hLYKhrkTEYyw2PkTaSt9cPzzYLpoQtS82Gbjf7AIVc0Lo7AYOUey7QyHNQn2iCbO42vbidVZ
pGW/RtZAUCew5jJJ1H5Mvl2p6bHGrd8OusVDBQnZlAuAwIGG4mSqeddy0SEBYBA3q4YkYcUlI1y5
zYaZAO4Ea24a92omumqRydPs/SzC8O/ZmqmcRWbHlPPZSzkcafFOcAMA81PFyxHXCJHRqBVpMSV1
6IWMkauMUq2S1YNyFwe8QhE5ft9t1qwY/upFxP1HjeiXzfV7CtTZszfaSlwZk1LNFe1ksa5840gI
zIB3R3O/I12Xr5fx8G1AaqA4MZL5bSeAnY0CI1ohCNN42olhX3aebiCzx1pyj1MPcOL4mZFTI3VD
eK08dvJZbjIl3Su6R3R7pfU7lpVoFbotebRyTjqCnKLyx3S2tIbV/5qGFrKEqv7auFs0zPQW8bbn
S4jG3ATY7N/5IGeB3TH4tV62RKGX1BT9LD5aslymv85l2WxzRH+nT94VjbAqGd7+gTbb2Hp4w06b
aSG6e+lxslhNPhlF+ezP7vqgUDO6tOSZt7TtwWKT5LJcD68CiVrHScs4r+bGdauIAVwZOBhvM1XH
r8IL/+CJLwO5ywt1bjdCEB/2Tjqnr2Ej6DzJxCjLZ5PNj/xRxV23l59tYLvwEs1e+b78UVL9DkrL
0x535Wjk6EkppW/UVVmT/ET8RLBNO9rsV0AizP5H7+aQ0mHMc21BnaOs+5RsxLq8uAbyh6A5EEz/
r319apm6H2GaUWCwZqZxSjvAPofkQEAuco8k4N/P9COhlKqxtKGUJGgpC5ndKTZrMuzHX14Stva0
X03OFWLAO6a8oTNms5r4bVkYk4RRvdcuUpn5PBrE/brXL8kftmmK/IsaJNEikL1XG/MZSXqd3RpO
EhCWAWW4Qf/cl4Vm4GLVTyFJ4WCLP6FzvJKrqPrr6/4/10q0QRPriVAvsLGRCjFXw51894/C24qK
hS0dZ1sFXAcDoQyM7fZ4Sp8BzYnS5W6DFmzdC9yIG7Dgy5JiZai0lXC+1LnWeapyfKfG0pZEERpu
58cgqgchrCta+d0ackO+JITTySESwIDDTbhjehdblCDRqYjjkGRM7mZOKElkoX5k0RTQXRiHnsS9
oLGpUikGpulUaPMCwZBNgU/h0eywModZUPQKCrFiiHArKpUDpfPMAiJbvTnAWpnvhSCFgiE3YQ8t
lLbLdJEqeRxam2N+aB7NRfQZTs8eDm03Qy5WRQQcypsJHhLbYUo3r7PpGifGxBuiCdScWTkik/ED
PwNf4Cmu3PTeKaHa/vjMmiSaQaLZRLOrwuDCDR0LPblUCJCFD/TQ2jEbOlqLRRH3dNOuIha9jKIb
nlWs0mU85dW0N4VIRHi+6RP+Y6D5vbx+x04hUtVuiajcmKur2/q7ZJUDZjxMacMo08LWDaB52Gg+
3mTb4rf60HqVHBrKe1WTwMrb1bSuDQ7GFRMaBhLdoYczG8QNaJObeEqkpua/OirFy0Fw3fbHSIeU
MNLGhzNkGv6b3/bblNgUuoKWZE7tRkQdBRoQuYrXOtCxQcrQ4zqSn6sHNPGjRXE3PxaRHwJ4QBEo
8oSlQ+PTTMC/WsokwCDNukbplhEJTotTym0NA64P96lZgrLlFxNQ8pMeuWVK8DIMeHN7Ab2/xxo4
LXvcTeEiNfxND2ubhFLh3TBiauhAdh7OfbzeXZNSTwLa/o90MRsCzV9EFPJ+ZDk6iZYtljnonlMa
tMx+6WWaOUYNDPQs97vz9+WCoriyB7WasB+MWDQvO3+SD8l3ezykpXzORFy+hfuufBpZl1kn3Hli
mZajMA/Jz+5XdyaDRfdFXeaMEPubBGIVh+O++gVA4d5DlFj/VK1A5y/reikkeHdXCntX0JEghezg
rwyQhj7CJ2S9jDBaTIFKc+pAZrG/6tifnIXSCWtXfwDrBGG0tfDiZxGr7YHbtpOTOkp28qatpDib
GAeQ4mIHyIvCnc/e8MMW1w7kK7L22ANpOVqQRGziLY0LzgldCx5cMm8Nu1ioTmX4EHCIaCwzz8W9
xA41MOSLU350AUCedU9HjsNaSzP7XAnge4zscdGOwwnwPpUDdeIzsVha7FuWom25tBha515d6u6g
UEGpS0lnQ/oKVRJNdgtMmKU2qi2bt1HCmNnHm3+haEEyotb9vWgccc8xTUQeUKci9pgDZm+U7+AT
kGT3YsLkq3JVo/Qtw76Vnz1PiPNypZdWLEqWR/+uy/MXJ4i6WxAFB61nbkN09lEZGqZj46jeSmzU
TzgYspx5Cj/C0MH255SwbuRC7lY+7v5wWVRgjd4acTGza3xdjAV5imVo0ZjDW0s5lFG1bzZF+5sV
NQTOiGLeTuTnuqyqyf0ed9XTg5NlEk5TGgeemFuQpkNd0KazDs6z4wyMZMz09K3l21GMa3gUb01o
wk044j4GdqUvX04EVNVqdjeSSULLqlsLmQbwRAJiQNQiGM05QKpCh4FBlKnKryqLNWNg1VMhbDiL
Luuxtw19DLFHSHM+B7SaAKsGexJ4VVVebF0Z0jnDc49CU9yePfrKUkEfxS4+omLjZsto2IaQFHEt
pumx3LhGGkeB3E9T82GUEWBIrwX6AKv9SpBWbSS2yR32v3HGU5YJ0P1//uFGuNIWX/x9a9aijaZe
RJfOCry5sqFsWWr/Vu4fYj+Krk5iUUZNO2PUhXigmWt/SJrt3RcCpCSneM58v27uFTf8mTtRt9yI
ufvtLMcnAC7tKuNEoARr0xnFALFIobL9b8oXR/Q/gyQlNZI+iuLiKDorlWnttH9RcvUe509e3QXB
lLL7EPw689nRMzpqA0BiUwUErIiOAc091otnCLcj2LbClCSgHK+OVWZzz0jGb2d2f/1WBYoqiiYt
RzLgj+lYRlK6yjzBclH+aX9NouNIgoTtqOiC2QrecmcqgM/3naarQpceKmbNE1Xv4AeRpfQPmSZh
DI8ABB60QKz47bjj/mMGzAWu8w6cQju00nF3JBvYNIZyZw09htkgBJkt/kd3RZeObjs4zXSNNEEI
ljdV4EVJeaWtI8TZogaeK0USgCb/AQuzoZ/3kykFtjMuePXMk3NeAM6wRUCdvj16EhzijxKlkmg/
wiGMhotg7KTeWXR3RHYODbIGKsg0Lugv8hYOlODF5oSWbsWbxudrkVBYRaIJw22aqkz6cSYjNdfE
YD1bbga1TtfdmP9+RwdJktq/a84fQggZUxXKPxlmEepEQa387flNv9WPD8L+oNMmNaH/ofgEHvTl
/zN1xxotgy/9aHWfmcdlyEJ+6k+bBXd1jPaKIaK/8u03+B667nIdoqrLgdMGV7FAmIO7+Ggub32P
t6uDd66EVg86ADHKyuYjzrFCS6z8Mdc2cJMrnfi4PM606baFOfLBLxkHRTQK43LCnm0rcTH1QEnt
Qyyjal2EsLXeq9DreByyI6jnUrqoVinuYzWgM0oHfq/lJw5Gz6pJ9yksjOicgabXBbH8fNm034pP
35p9rmBEqf+lWDoU4krLywL6NwS/U8v/iOLQ019GLImpSBkyh6TlcgOmhnPSXTQb65A6/Ov9pkDR
BJ57V5lkSKZrLxkOI66Xa+m3edvqM9TDaF5fE4mK22geyraj2CWhh28kmwH1dz7tKJ24Ee4dwD8f
9M/11wVkF4bvFI51JzYLhuuXOOpqdmbuq7O60IVzFGHevd1QOEhkTvWTUXpGPRa6SjFIcdRtH4tn
Zs6PIgn2S7b6oDPBN98jFcIKVkPKFOzQz+9dgL2+L43HAqghyPPEItjcnoUmsGMta6U0PplGruYX
+JXpiQFfx1nCUxBzKnEydo8TLjQlD/WeZ/UqHJdt9Aqgeuh/Edy1P3u+DwgRa2g2R9gSx6FAR+Rj
dT3NUS5n7+Q2cpvXgpfanIBdVi1Laz6KVfsFChLS5L/oViSVB0lQ+YSMdy48lQJGZZlYj7gprFIl
sGONhqCYsvNO9FrHiBs6fvHhRZwzKuLyfjF3z5tSsRoiM39hbFw1/ggLJJSnG1O/twEXjxtVbLuR
jPKS8OZniPfwebpBHthQWKo+bF4h/yymqJQzsFczk7FZk620/JcwCrPJxTapVjaIFOrhCz5ZWl59
wztGo2s+fP0TmaInO7L7lLzZWRI6/OioyryV+30Hz5tWcXrtdp6Y8qdkzq9kmuKYPmK2Lt8P5tVh
GH8IDXiuukPYI1Pt06m19YUlG0Kw1KQ/jT/v18+V/xzAbzWL+iALVB1MUrPbHgpb4XpBtYX55ReM
b0tdayla76wwU/n1rg39z/uFkReHYokuQNaJErdXdLT6aEKO83c9q9atrd5bgzCuB46Y8tunn7tu
rT8agdx2rVP6jAMsw5TCmT8RDVYMOKrQ2ALUE5dFlXCDqKcnSzMydmp0dkUOtgIcovxFKjslBJ7h
E/KF64RJ2ZTXNX5PdKiGikhHnXt2rBFGFvA3c1+wb6cs2bz/qNcFCcv5Fg/rJFBvGRETISHMKcyI
W5kCB7SsEdL1H5F2mpzeOcN/pQzonuXp0njD7rQqpHydpSKS8HgltcApWBLhTFRXCEdxNdzidJ+i
IsN1I1p93Cp1kASefG2xn8qJnXKDgCB7z5N5N0Kl45vcpGFMwPJvBxxCMCYuE3k7PodrlKtcjvcZ
JRATyFOjdQ27kThgfZP5PvSOZlZlPvZXQzsqtJi13oit+CcEVrdl+i4UzPbMVIVDKU9E5Dl4+uXE
7I/MP13KSz6f2te12P5cA16WeQnq92440keSVogODRf7kFVF7Atf+A79esRw1GV7y9MmgEFU6wDD
IMtHB2BnRWYp43LgWyHBZzRk6iCAaYHYulnekicslWCe7m3e2NSPjAiZu2WmgW4Luokulmn6gUVa
pa1QHABHJQ9dUAr5lGcnuN/hAyCeUIuSJe+/FHusSaKqkO0SFpV0EqKNN16S5AP10vDhmL+CxKEZ
B/IaJiqxaZN+YpOzzOGGoaxrZlUvnxB8Re68e18MIB3FmyV+yPKHVsEnNNmqLw37HbKA4YFTjyhS
D1Htvx13kY/aKEv7yZWNu9G1N6dU4HAV3Aj3MWyBDGlDylDg7bKLbHNY/pYToG1rWSG6G7Qo8U3g
qBeFMIx0/UDg9tAVexGTgNemXtwP03wb3LDyosxPpJqMRS5pI8oDbH2oZBLDHjIJM7v/0sWBQhrR
kBqD31j15SGSAlNQyfmaYSpT6FuzKAAqXCdv1dm8WbfYCOQgRaUzHkbC7Q5SEYvUQsP8nT5iVmOE
C+vGreCsfuT7odt+9VkOmRWWEFb3Hnzjiq8br71t6ccoYa7VPXbyvXj/B3AKQE+AqwEckCVuMFSM
JopmxoMqUb88e7tzou3iq4i0fUFJSNAVwu5dVh0uLCovTfh2Vovo+Qr9dMwYHvt97nkwJ1Mz0XiD
H86snHyZQCQQLaHqM+pJOSfvH6Xoc6DzsTGUiJGONcDXwzSMs7pp49DlxhL+0nzBtXwrYi4eVkhI
g9e5pVferw1mJvw1g33yAv9FOMQ4WFqoi7vFKTOxtDgxby+jFYigH9bR5wGHqR+T2ujM8KeImW+d
OuSBWBcQBwDylaHVAC0BAwPGEYbQSdwZis9udkwD8mOf4l5BchyuEm9DmBojwZgE8oZEgG3ncFls
YRjgVeskKHrTBwW2Nkbx1aex0VhHSwaK+8U4peT7iRIq0lXowNeH8ETFbCo4fX8xeiRqh8Tl8F5M
MJkUbhk+fpnZe9bAYO8CGNqpSLFYpZwtBt02lBj6cUVtOB0wt2MWiTw6dZuVFigVTbxVCNZLGrfM
Z58RD4UJ30ZBU9uJa8WiqW+BCvPAYsHc+RxRiMjVXs25EatkOj1Yyu/wdwisRvPb+7d6nw3F1C9k
CSDHXzZwmlTZviDSVd/qkrQ27m1WAH5Qi64bGL7ZX9Ub9dpHnl2T6CYXbvQZKqZKn9dvhkIT7wk/
f5kSsc8Q+jtoQbfWTuFfR8GzMSL9nF6XNWMAxPy2kYJthY7pUT3hM73DBqXbPxfVYlqjdtEepA7p
l8dw6QTbMw+jRnpY8AyTI4j/sfsOIKDnAjAEFzO+uI+XuGxRwxeDgZiluJp7ZJaKB5xlzKEb1qZu
KuXkT8C7sjLeEmx3f4V+aTNg8LrX6zpl4TX2b9SY49nHhEAddz8vkbJW8vgaCJ6ZfzGlkAIDZvDD
znZovK5TgzP2bhr6YURK2CgpB66AGJDUU10tOA49IdJffk6BT/DE29v8gJU0xrI+ES8ZsNcZqtYD
yV/q0c3vDZk94SWQBGCEjNfvJzCOzBUCQ64Jqa5gKOlIRDR4pRb+plhj/gLeMvGgUoR4syExx/hl
r+xU04BVQAF5mIFkBOf8fCQtmClTpH1j24W/NVFDJYiQuhKWGKLGWZwUt7i9j+CfI14kC0+run6D
kCq4MPwML10nHeQsHxS+/I24Kio9F6XkKMZPoAYqON3iRdwfGOs64TFjCfroDi1lDDC00MwS7fhE
UuJ6893uY51wngihhY0DH+Lta3dSu6sE5RslkpCzT2e+aXei4BBeUHtlUFOyourwzYSe87fFx529
kspWxY1uVymTfetJI/w58GCmVH7uDMglL6ssV8q+7g3NN5lm4Sg7QcvOysDzlwzZK+kWPUc0FyJp
3Sd/IxIR7idjv18tPW0A9YZX1XD7E+2dWB0CdZpaQWCXPKw1OXKBWsjZjYql4Bbc0nQNAaOuguJx
zFItsGEnyhHX2y7mGguqwlOhYArBps50C5gH+ws4BEcYAbUhmlUr1hMtlmziSZF4WBtOgS7Ng3Qf
N8gBuX2qD+d7h3KFOfTjrOfatgoisRSI/ADkkaz6kiK3dl5SpE/GMCIsDOGiESab4h736pkpRfmk
c9CQCavEWT4y8f1afGFxMXRBvHCh+zBnsNMQ34g3T2IX5iMr1050vNZWHcoTy6wB153M6XHtnHNG
SBNCe5b02XOV2l4tiVqos/AdJjBqHof2OvV54DplKDb5vJpUmVmHirGtDGIIjZPl9NDGJ5pN9D/g
vFa/IUznanitaK0LVXk1hRBuMOxyyyyFvB5q/7sOw1i6xbL7eszXTsoTkubV9WjPhgdTzBTZenAI
tXFqAGdD18JJCHTW+rqlKpJlQNBGIiXOIwU9tFz4+GoOIFcjUaApVZesDyraBYLJUvCAabPgSq2I
Vi5KeWYo0p3IdskBp33+Ik7nD4Bw8J1snJ1qfgvl9taA5CdxSG+Mq1iHNubEYDij6d4T2y1UV3LD
7WUhx66YDRkrZhNuQTqtNOqt5nUuc+fTDQTPzyu3B5yZYsu6vLOQPgWd+5a8iJk+puw5bALM3lt6
hCPUSgtn7BFY9T9ZXU6A5WpdAUpDS+7czF3PrDSdfe8wXq3Da4HMA0n9xpVdQb1xhG/FGjsNX/gv
D441vD6n/ISAjM8ouhQA8Lemgdox615GtaPSAp4DOFfGlAcClsC4F2q5MwmMJuaAbGInurmNYOHC
aPld93KivoN0C1wAKvDZL+PBQvfTNze8iapW7uFGEi1rCPgRnokdTlbPCOaeWz6VQKQ2o1u3Yp/Y
V6s99UR0jENeNnALVHqEHmGMc6rOagkZx9+SVqQiT7USdOyIsxMbtrqBLqUv3ywbQIw2XYceRbYf
WBp4bIcLAWRKrgqB6tpdCry7zXEUeMqa3O/vVixwcRecOXWJitXtr7nFopX22XYL0pAZKC8ki2Aw
8bwDbdqp/OyOjh5/z9Za1uT1fYTDxWkQb9EC9RU3q8fpCCsUPfhHAGRIsEnmWsChz+BY/8WCM+kR
SXyS/oEIhqsg//q2IVso5TKIx6VTkFb8kCxoMHdX3wsde2LgY4HQNhWgSHfd7TKZiTpQL7jYegku
oiBvclvcNcUrK1sUIovwEKq7PkEq4t1ImtP9U0mnVuNQS2s0RjOM3pwUzgB07Pp17Xnc706o3fVv
MRgPPL9/2uU6HXP9pG/3cYGYFIusPr2Ph21LWTgJMvDaWqmoH72UuRoYVAkiHDLII+F8HwI3LnXz
HT39bsGYGMdCmPmrgm7vIl94gTW5Zxpd3sNmOocDP94YyKcQHRaxqi3fh1EwVzMNSdouvMuwt6fs
4BHjxxvCOjyE1/C4uzZrVfd+tsZ52l0bT6UQk5nwhitje9YQ2cgWn1t0QPin1W0T1eiKasQyUPXA
8hrjIedot6erkpeY947c4x7MrWMGmBVAQ+BKP5C23t9/2VTM6Z7SR8P9vxyFZBzRiuu0r/KWsdFu
RwQMOJHSbWY05lO93mM31Ms1Xld/ExUCMWkRfx8Q79vqh3ZAIfBc0HtzDfI8pTybS/EcnYy3Ko9Q
oTiBBALhl4pZkPFjONaunyku8SyKuN21aY+yAZZ1bnKAuCg777cqUkOAYIX94uIWY53cD53dkYdo
Y1+XBBjrudFlbb1zWMbPOnnPOVGeee0qtlsv6W4hsMEJhq9KdZ+BDC2r9EbeQmHWToxpSlm3i5oV
Tbu0s74LKM+uPiRpPRkRutvAcjm9OA6eP8cb+tEZF+1JjdZdIR/dBSxC3O6A9LVgyfPLLeMFAU7X
2QUI5mDutBgMzHvuqMQxACe42ReSTR8GH6zDJ2AOWJNWB/nfedYiSIGiaWgaSm/P+SO0rqhQeAC1
tsdZOrkXDRAx1fwfWrerjHSw7erPtnnXCs48F7EmzVujzgLhw3neObGnjkEwb0x4mwu/IUPjy6jX
PYru2PowqrToGgvly5gtfKfVgBgPDq2fZepvAj6PJ4L/zw4aK1ftiBbm8py6et4/Sa8GM5aNkWQY
UYoamn3WP/v2ngO7a+Dqrjj2FRqOjIXxx6t92y5BFwwc77avmp9d/ssOocWCd4bHuZuKGo8ybc7u
ClD/x2eyvd9wnZL1dY4+mFUuSDGGLrLcdJ0UI+IG47RHPYEqYdX6+LAwl3nHTwipvfqAvJkBNyrV
rybRsw/MOhtN2yv4IaMNwQWx9TTd4strBTeSqSGlvlTiq7NTN+c3l7D5+jFjcUwOx3WPkp9LgIux
gz3G64NcKj+IiDNSHrZGXVLiOUzq+qVH55+Go6DcxG7e1SJOUsV070bmtB9W0Bk8E2v1HElJ6yIC
fc4IctJfHEjZlhS+RxpbbhSBgtIv6hJta470p+yQAnvslr9YnWiBdxXZvkW2H0313cbk/cWAdTwy
WQkqKZ30/HwAA5bOzsN9iy3v85wEWjJ7AKRmbDeSLUNb7/6uu38Dr+tqgdOhXybsQPfaSrs/ASE+
UEPkHwzjaAEiB5q2ZI6XKTRjApGkqKl9GDQvg+RVYQUxOIx5I/qlmXZpNyLan+XXQuQby+MYGB6e
8O3Ta1RHLjaP3oTyWad9iCebdQwxflY++intS+rMT3vqaRfJ462aqLW73NNuhD8+FT8P6FO2vbpk
9ZXIc/Cd1DeFmvqwPVujm5JwbpqtURusNQ+HLZx2DZit4eLcxzVxgXraVJXNGzVenjdd2RIZrvG7
2U8aP2cmB3HSFp2Wv1H/PtXJixsVWrdOsY/lsNph/we5aJyj0ZTXpll+ZOmkIzz5pUr6MtERVxlj
fZhJubfybyhjvK1OiJcWBjlMKfYxUkJtzMa5teSn+XtON5CNfJb7N/bOL6VqVvsKyvC+81vZYpaf
gV+Et/UqY33o6mOTinRkzEM0jzfVpy83Am1T8GGjKdhh9idZCcffbn3aIBQpiciiMMWap0YpTxG0
EJXccJIRFkHwt/EoVmXBHZ8C19nPqXQEqGkw5oWzp1lJ/FugipA5b2XMeq1KmW0D3vln/FB127Uz
K6FKmwlK1dzdeXr8tX89Nnvg7LgaLilTfv8bY8rRfUCF6WW9YShNbwV2UiSRyVbuK+iTQtFwOYxv
VIOWvUmS/4jM6xdm458wKFTJPlYPbMh5QLbmdAQm1mQsfkpRDT3+eqDjd++88uQv/vxPwangulNx
+zJkR2yL7UCvMfmzCk2NOj2ycHDiejjVmmIJVlEWjpkXi8yIeYZsPz7Cd8Vn4ILB707PATEoAiHt
sdSgQXY/pHU5Kvtr8+Q14avavhnlbvjfrmMdvExKW40z1EtivOdG5eJtAm2z2qXZyIoGd0PFl1QD
XEyWOrklxIsl62d1Af0DPjd/rT022F4tNExiw65TQf7m2O3TrD7q2+a+v1cDjLQKxkp46eUItPlO
phF5VRdow+bBhGPDAnVmW6vnphLS0N8Mr6qapwjOA+NYRJpELcefbVuUi5ED2dHcQhw60qw3n0Pv
87mlSo20Rumw+zIDnNuwY9m/klbAU6crc4p43EfBr+TDCiPOI0+BjdvNglICiw9MypLcxWG0SMdw
3u+6e7/BVdHwUHCWszlLydzWQZ4zcDz31OiFaRkYlZRuVDYzG5RD+1YcAY5SwmZjMk1or/a29hP0
wio+ZED9B5uzPhJ90NIeHPqI3HZKBpJ4Iu0E7noegK1Eq2jtXYhv095ZcZ1xa0JVEGAvtWQCluY2
R8SCpxE9WF97l/iqfDi19ij3F3RofVW0qi41hSgP0sDoLfAMaQiWzL4IxSDL0jOdeIppqzarxHLQ
gjK4rscALPTQGC1o8LIglJALUKZjfrX414dAPQuwzIaH8ctX33AKnh9S0heW20h8dNVbHhNZ6pbh
XEsskM3OYCVYmAkXCX9S/oCSXXxP9Y4dksB+621OfP9ZZouoTkF1o9qdR67ik/5xefuZx07/bSJz
s/7JJHs3agAuqxA84J7/a/TNN3Zt8FXRlqABoVksNwWLrcM/cRuLswSePT6SfFqIHrTUnP8qbzrf
InF5D9/2jlbMQMjLeT22pcDDPwfiP5hDQJGpQosqbmZphV+WQ/EErMikzvDWQoJk0kX9VDn578aB
KBa8yTyasa2Kx8+Zqfz16L8BuAX12jOceTF2l2YoQClU5wM9GMqBooI44dHEadgZpi00GD+a/N8R
7UYmCibLxuQb/fYF8/oNxMSa3B/rdiaMFQNAi7ZsJ0n5FWZdtpg67ZLZaNEiJQmYeUu3XDzp+Cuu
KauS0LpgSZtLmNd3hcr0k3yWm7+C7V+OaQMosL7+bUaLX3fRC5GLW0OSg89LYPROscBfT2zBENAE
SkBcn4cVospNxfnU9BmOH6Z7R0eWajcwVOkmSe1VGZ9Zc/K4cJ/V82xbRGrFiWTB9JrgvForPJTY
a4a4iuGLQWsKdOhCXtESlegUMRVVKab8mnWX6x6mHuAUlpyjJMmD2bmvNSMyJBf4SNkA/9gmAV2o
PO3NQZJGfq+tnBY9xo8qeUaWh1nU7Uh9QDYku8RxZZflG5mrsY5qk5PuBWOCM73X05mVmDuq+7Cm
BuN1Y3JXNXirsfBnecv9HHYFfum6SDsUbHgN8UHHPOY/ZfbQ32pNTfDV3tcOD+5r5EJRMsvgQz0P
BHb7cS4OMqAkPDIBweJa6QO3xAmf9SzQfJdXf9E54EchxmlUpWSYBJ3GYr+d0FyH5smIKsiTJHa/
EHdzs3JCH41luwvEKs44rS0xED4SroofvMbo7CpTZqBz0QIYwCeB5/jfNG3CnqHe3X0bBIKIfUU+
ZxL3AHd9H8MkqRI+FM19O+mMQLqWn7OwVRRWyXb4xd2Xf8/1DZyzBp0OG8r0FSQYNe4ZDKKSSN3g
SOLk8m8IByJkD/KxGF2Yj1o9dFRq7i1RNy4x0zjiMa1D25sB8d1hFUqvSOEOrQ4YnB8MzyJA4XKq
o9KQKWcE4VmAXBZpy2NiXJEBi39t3OalX3rFb0mgsLsEk9OFxlMwHcLJF5mItPc2GVV7aG5OMLrK
NDBCr8IPDo1sZ87FJIB06FInyJtPIkCUCutiMcSbS5JuURCmAIE3zk0SmMaqwGLLYwOm2YLdDH/j
rS/5lXvvxW1pTKYhXkWKofbTgkuOpTspH/sdBPTfG4sAtazMpuLWjl6uYJHz6sDIdrMdWgYRI+9y
46wfYu8ywR4TtQ7D6uNA/DHauTZT53g8SY/M3tiSYuWk45d6qg71PImNpWve8S34qA38j2F72fv/
8Qn2XSjjOEdCIApXez3Pyqpen6PHgKqgdt2tIJOdfrg2G6B0GHjC/OFE8J1Z8F88dpaDER+v1O5J
qeEEFjS07Ui304tEjCM5/RLUu2MVC+oTpVGev7tLTQjOkBQqTF1vdt+U5rlzsyv+zmjpGsycD3DX
uP+VaVeLjEHvVxdvqRLkNVoNyAOqjWPwVb8VhMZGn2p7Hl8T8W7tyDkEUfqibzIoIlPhQc0+Tjtc
jhoKsvYpxfSDDdaohivkULZofmVvayfm3Ql4zb9qhnQLnnKYQOXmUl5VNIP/F8u6izXx8rf2QaMj
GmM4K6kjlcNbffa9/s2iS3jAFH5Pg5rYaABjsoFSnHKDMwV9DxOyDFOuBWw+T4ugUFmy/HQmdrpr
AeR9pJMWPrjmTEP+xfhBuy0sQp2MPPGqfTKkqQtc18HlhRZs6IFnWB7dNwWuwqR0U49T+CtGVW6x
Xs0Td7tZ5cF7NIPkV4Lc/YdQWsEqiBjlvb+a3E8x5N+iljANBiQfbdJt3fT9++jhY5yyAlgK4CEL
7PXHkodAAu3/BBOHsA32cHeqnHqOLBzfKzzILSSJQSqZGpGrc0DZhM0yGEayn2aVXGOlIkapgKMR
gCxxYXpgn3csmLkYV4eG0HL9mtWTLm0NiS14+wrJ9VJp9UJzeftd1cNE7MPZdbzTnIR1EEe517/q
EwEK5djYznOW987gHaQ1ZhiIyoRKoHV+lrA0VpZVc1P3LbIzrNDvhT6Du8UIv/ZAfeB+VV0IObkf
XaIW41ZYFEkHFqqmnT/zDW9Wrqb+kOZYWIQx4yI5kKVWaXJtxyvoCZglcHK0ndDJkPjGCU7F93Wc
CFA1Tr/B4vQk2wIN0SSSeIj06dsr/CmU+kwisjO66/qeyTjU6P0TMNaKOHiIiUC51TYvQALvNHkZ
OS9fr7rz7idBsqdnpXpdEcs2TA8VwonoeHkljUPwhwHTDJt/v7aFdMZuYxOyUmWQ4L4sGqOutNr9
lOhMa3hkvohfrlNDj4gu/vNmKdqGHmDnQbXJQb+SwFLt6hcEzMk6m8Utz4ld3Oq7WT3EsHPV01K6
hYVE2m94ucGTxVVsIg2IcjfVBXFnpJWZGGl9Nv06TMxzDQiCCvEEU/PMa9c8o2GdSPh4mmZajFve
zyVou7i1gDbSyCqsm2yfWhsuv4v96OZsClpgGw4dEAhHJD9qTz/gIaKBA95p85mMfrZvcRdVBHx5
AvDd8Ub+YF18s7yAEckGDfvpmAPh0iRBfDmPMNI7yryJamk9m4Qmzi8Y+i281qpPKF81/3jiheYe
GERX4qqPIKZZ+kkeHqgSM/LkbyrXSXYRKaBuIMwZBiH9oKQHDiIPQzr6I712VuWc1Hj2kJuCTHPJ
U/KH8nPqH1sxjehmOAx0Ji3u/zHQWh+oz3f5APqRAnaPOvX2ARF+Ml0edy8SGV1cmjSbbDWPoECZ
Xz9l+H310SxKYc1IhURZtwRx5LlMjaBmt+7uhnW0cZINq+xhLWslvEMBldB9ifIE7L6gdqMJobRR
lQ9yLAwg3C8YTDH+yUIPVILA8hBW4IwT3+iYZjwsAxl5pukGBAuz998vncH+Jqz8ombPpTokB6ih
v9JGzohoNAfbu8KMAHcTQ2zeHXrGAEnxEtJZu7Cv/pTgLar0EQ+GVekHZaDiJqRtSH3YgWROnDtJ
2BSXUKMgf2IYGOV9Ce2yfRNIWjZkRQzTA6S+esx8wKu8eriBfqFJ9bJvcpoXMuL0riJuUfarX2KP
eFX6TeH+TiZGecmBqQ/EmDSBnoqNDfRU9Bjz+yBTmeJ+Kh6JFS46bz72EPiV1HxW6GjAYIhTT4gD
mY7Cq3fqGnI0HQZf4frKAYCYDNbuok05HrdmUfhrCZFKunvfM26itqYWbjKTjYmY3mHGigR9yjG2
sC5vBJT/x9sfqWhMeLr9Jpy7seQimR1UH/iQXvti08njYg76ye0sVpqPPzJTh1jdPbMibT+wgYKn
Alp7L77ZNXJY4dzZFaLMoTYOMfRQpot3PXv8oRjyB2KLxW4ccwdz9+2MgcZv39zLgD2QqO38Jv/P
ZY/dob6AEFRxJafCKeLnS+1uQp0Homhb9RwKNkapBjrMowIzUHBTRzqwfZ7wKfTcXaAWxeXXrCqy
8kErZo6tVOrulyCWuBu9YHanzEGZ5kO7ycAB6BGV1WohxkxAynrnPOUu7pifmQQ0ACXwy1z9xdfo
KP+OgKHzf6Ej2pqyxGFX7fCEKt7gyrLm+VDueUPExgRPrNkiTV9FqOKK+fGkiZkSOeePD2rBGFNr
y1O+5xENJlkxesTbAINB052Br7gL1iSI0WTSxhIqoVD+tPDoB9zjVf+AUI3oAgKjANzrFFnIsV2F
rkQ/AqW8QeCI4aZm+otqDlZWQneW32EMm36pa5IzpJaJwah5T+pKBEoagpFI3IXjr1wFUFXoTA9k
/MidVUqwept6sAq+gkl7NcdGVHcUrs6BqtdeeBeivNEkohjiCsRLXgeRBVmNBaM2JaEJ38UygdDT
R5i4wsuCrTl8WLtZp5dVkA1Zru4zmHV8NmCQuhKW7k2L3QcUUTg6YYUrn7BpXd0CFRf27B75hc3t
aHLrypBtPfbYdkWtATDv+nKiTPuHYlV5rjYEZSGFsdqk/iehoZTSp25olfn8wgklDGAJtiwz7ZVv
Tp8KiTS4aCocYQui2EKgppTZsCkirXVx6kuHDMzswzwVU+lYVVaHnXpobm+7hItgUBYRj67cpreC
hJ/q8J0O89I6a2LDTal+U71JHZYzZroYCqCmxy2iRqCLNmvrXB+Plx6tkL7ciZI4jL68JCpi2Qpz
ftLSt1k7knIBcxv4sAXZzGdRRh2quxiHy+HrMx9Lccd8pzmwlsCOsQOJ0Rzv33UsLLuvW6WO5q5r
EyvBOuuGIUzwM7/SjaDDtVSxramUSV2o1ytDq8WCJCGVfQacAvUYPPpVFKRolX/C5mCX8Q5Qirf+
MFBcps8Iil4g/N64LgWwvgd1R7CzdA12ycMZQxQHenOthrOd0fcMV64QWSgkBCxn8r+NWN+OKTRF
B6Niv2NNsacN1KQDQyD5ibO71UPLftFAUs2QOjUN+LxbaeYsZ8N54zX5wbfxORmOPGBKdJNd5hMH
e+WplFUlmqBXmFGzzVpLnvH6qrm62bBrxCVcKcEvRqyABljnIgOugjj4NRWv0RHfEEe0JXw1oRlW
y5SLlOqNSk8pe5esUZgm7vlZ+tuXyKipSfQHbWNhyveqbpARgfz1rCQEJUbd5pqKyN/iUnZ2BIu3
qfNY6sIcNT0lv3JCyZ6jlbbnmJhKnQUYankHHa4oA8xj/UWZTOuPcrWWlxpqJ8nMnkj+r9lPLXka
nphJesCrxAOX4nQT2l9ellzRhZBhgvXkdfyhS60/deunlis8RFIk+trrlJap9TvRU8NPIyDr4POK
5iqbKLahWcT8VZyujQOipQM1M8TThj9tZG63YNS89PKm8xu0hdmS1dL8vrT9ZrNC3BBZbsTt/li/
o/Tmj99Mr3rgPbcewD0rqPjD/N1YciwcrxI5aoCXgB6iuMc/rhEtQ4pm4RLq6s0ge6YhefgYAY58
XOybghCjoa/Fk7ZRbyNfVDoteVhcP3mikF/zSiF3CPfF91FyS3FetT1xvivNpwZosRXrpt3PF7Aa
RoLlNC/I4FoN5e6FgAIOPQ11ZcEwqSHzKMlfPzzPvit0xOsvlv4Hp43upo3Xm4J2GuZk6CQQKOkj
6bzGiPfiqwSUkbFAINnoNuYHNUn/GpSnrkeehHD3xoovl/WkONKjlsBSIjB/oPKYk92d46WwRuuZ
caQYnLcE7v1z0u3W5h5ZUNBBvc8fH1OsnhiqpZlvRwXjLJW2t5ncG/Pjp3FB31H4LA0CUlLVNAH7
JqXWyN8ezEmmgM0X5IHSHFPqRaqIA9I3kvBWJZh3eHmGKqKep/Am17yUIZdTl6b8GA4y7VfhGPxe
Vvf9OQ+U5Nn6O4BFyyG8Iq/Z0WJe3VQbaHxgalCYH+QZVApjnVvXa2ggjbaQhj5zHxW9+aQ2U//p
8gSO1ow7E0oWKrt4pI9xdBZdzjWfzf8O3DQCxy7FxOkOMhVE/Nkb7X4br5b+BSEDfPsDxcUP6GVa
xmfLcMJNULNDF0UMW7Gh4UfhIRnO8pODm7dy7IpIe5X0Zufjji6u+ulbg9K/Xf5+dpAH+TMF6ddQ
1eqhJqhvvfoFMwnd+Kr8TAZl7pHmzyI1vvXKqiRwauv81Wy1qRcMDS4AbXIlPR0C5EBfTNnFFxTK
YjRpJw0xElZRudi5zcYwOYl8SNfVRIJMLqc6pHbopZI7oA+UsDQ48M939/L4ARxcp0xvKBZkMWRI
N7oTigZUp8Wau1+lxXzpMKY/wB6ZPmwBvw1iIqhPhor+cEMF9XvFNX9P7oflICC7Q1vfMhcNJdIk
sXdgf3p0tAlIKYLBpk56b0SZuor9n1+QTTzKg0D8KMINDtQQ9qS4a4O0M/Oj+L+/C+kGiZ3zFqIK
v1tWKExfRbNUcXZeRCb74z+er9fD5WMnEntN/aIJ+WS3qzWSan/hBYdowuKiQ8Furz0OSq9Cv8np
OQUJgjDZU620MAAGALzBgemTaMZEp2T+q7V0aUofXo9eFC6uyaMiCmynvA5Q2woKtm/2teQ212NM
CLmUH1tWH+CLWsUw+FV2FUTv6iWNfX3J6JMzc7U87to3+nm7zfmdMoLpneF0Cv3l6ULC29XHPdFV
H1oXSVKE5gkZm3XxZMhJ13BdmX/CA2PuIffvKfI2M/fJz0a4eAkGZnQphliCRRrYeVdSKjLwGZOl
34U/p8ObNT4TxRIyazx9eHwKXwuem9uUElyDUrXVEK7e5AaTKh2M5RqZK86HfayykVr+IpsSFQju
rjpZBFy1smH5ZBZATLL6+oLSjSC0Jf4EA1NVIvwF516ttOvooW31lQE8HyJSrt82rz19XdzgSie6
U6WBiOaDdDiEXHTEQV0yc+uT4qG9TwhKXlVtdYFt6NKQsTu4qrGHw1AkfTIFT0hRXRWkwUngaLJm
A9JK+SWwKxz3owGcAzWDrlzJTksk5QtNSMyVRQULmMrNO0jhueY8S5PH1eULKEAS8YhBAHtXPVhh
dYtG8tBvpfo7iHLPgeKqCtyhD6Sjs/v8WIezaR605lsE3j/4uoewgtbl6CgJDJOvyO4qhi8Dfvy8
Ec19Kl2cpjFGfcPaYB2poMn1W0U9iJJkWUQA5YsrgO9g4vhwSRTd1LygHOG3viGL6ehieEgQuglN
xEU5SZMID/a3BmVdHxDyx0/f1TJ7P3Hyh9Mf3C0ZueRmdDhDfMt1G1mTD9PDJrwJYewxljNSDAQL
qkaQaXkflz3N15QmV6J/xhApnJao/yPOvL8MKxZ6Y/0gee7+28QrAEQWz18gpWzZMBJFzty/naA1
IXoLRoq2OajN2nPC705ORkGn39bqEe8LZcKN/89fVP3Zv0cERdXWCuP27aA6imNvjZm8DoRvAg5k
0+Tm8eS1DS1R4bzIoL77U0KePspwZ+e5ZK9tU9SG7DRoLwsJmrd39pQUVXSQirW4fDGhzLq95ujM
jUVCDXMcHPv93MtnvVu4MO8kX9ua8s0HqOytv/v/Rab/rlGTUwPINg/swfiK+gkaGQ/ko0NmhPtI
Tfa8VCNG93BMb4MUszJiXsgmmnsNoDGmX9Zv0gw3j5lS2P5KZStEH+BgolxafwKd0lPsDkQW046f
YphZYSOcZMVx/VAp0UGICRfS0ksaPYcG3EjQ3cUFmkzTeipMyJThjZBsGJNbc4fgVI5zBCKQCYTi
KEX8LxQifyPcpd6N41rbjPdGShs7sLPvvu/3rpTB64cEVCA6XtNSJc3zKl66ffem2GCowLcDmNba
V3UTI24DwJV4v1aONQutbD2qHZ4Ttwe+VyTiVpL2NTo0aamI49aP0PAv9gnk15BOZh42cMYNvLa9
wNskSk9AQ3+JgQlI9ryxGuMe9c4bBlz2cV7mPYJtV3/kXdHXmxu/xm/V89V1IX49VoJ0+6d9xh6I
mJiMSICIa5K18DR9KqO3O7CGkbH1Q0+DCyZJGcpS5IxDRQoqYzDUXFVYHPDM+Pd0DTZluwFoIJOA
ai9Pr07FzfQg6XZH+r7EMtWaouTJS3Ar7SFxnarOW/VFYGuYQ9ZM3sFePF2dDtmmk1IqxX2RRxli
x9/7Um4zB3doj6p492iQwvgbb16GxO9fKG309wVLgEKRV9HGgRma2O3n6yhxLz3xiptGCpBkS9u4
jUlT3/capyZ9njPuUegNaaOMGW1mZqvZQB/hL2TqdhCpA4GfD0k2Wfi97zT/w7iYeo4bSBFpseY+
EuffqLJOzIgTLTki5UUfDIvl8gim22QdjyZuajBnwlv8u6ft8TS8dpfGTNkHE7wuwaPWxbGSpKdE
yDp+ZkUXJbm7DL1n0Y4cD8MrXRHMFtLMIeArqGPaRalsQd3S1Je70/zh3KRH8p7zzQdHJ89xZHDW
EVP8Ori3NkU5mVmG9aSRQMWfxTfydWAfKB+xyYVKLgtD+fg49CkQd1POHJSNDditDItnWsXMfVRD
6fGMaAyt/PbhZbLUfLOUaY9VS3XtowcplGYxEpQ7I4iLyeDaPnpoH/gQOhzX2rXAtctrYSUpuEsg
SF/XYbRHKc4xD6zkhZNQFk7tqaxA8PP7kL69m4ohAkh74TwGLfFeM35NAtfQ1UJTKm7ejcs9cNRA
5yb2MeFd/GLYvg05dOMKqr3LolRUdHX1Oou/Qs6fmZQT7ZyBtCieXLI5gQ6oVXw8j0viAPab9CFM
2teeRYrapeLaFSq4KIfBGv82HfeGs29tWMQ9qTfDsSJqV9VkWhEH/5QUVV6jNrz/WQuSm/RvBgJW
X1Z/Sm5bF8nHSaAk5vrGVAopaSig0GJlI7JFmc5nslFQ5oz2Mw8rBwqASLHl5n+t1rpg8T87rtyQ
LCg14ZAgJ2JDPlLsX1JFka8eca2cjGTQV67yx31uI/gM7NGGxzUoJlL1/m3+WPbtOy83u4ZNS17p
i+DQvwBdeRhAJrCFg4OMAKM0H0w+zX3/VKhgZKJxBQcXXoFeOVnDb9Am47NOFqvJQbfiggQMkxVz
7h2/DbPny1odr6D2O++nzH9VieJd4/1lb+EQhtwmVzmv3fnImM4pA7LV9ireDz1Z4sDBsuB7KBQV
84reSCfQu6rSIVHNKkxLezXLx64YdV0DNTGYZss7phQ4XdiFNMRDrqqYd5WyxLDKnM9zdVLIFgRb
E1UdFqITN/HqmPdAsqzVW4xFAUfpk0VJGGjzQXZnnZzcm0MScbWkXVzjSlCuO+5SzvZCee/iXOda
ifD5iNVtLBM0l6o/tqVdBYXACeYQzjTeszuwRS92nxd55H+kDywrOHC5/HX+p6gTqO+SIWpte7g/
i2VLHq9/OlYwSunzfl6uV59q4aT0Kjewp64p4uCsvalcYaWK5GQvgvC2lbzNwVFdO74g7Iirshql
nDYvAgQWaFrdanxBfYCusqqtCPq6PIcRW8j1s17Ra5KKWE/hz/OrWwEH57eO1XRWO9YYV9ec8CQu
UIeM7C6rPsuIbly/U2NveWPG464OI4jyGMekegLVCHUQg6R2HHaLsul80bKZIiJq7agaU4U+B0i0
2oxb1WfoW6sI8xCkKdG7OzGxExYCedap1ufxdSFq/fjPqto75QqJPjA0IyrYQQeHlkoX0Fj6UXXe
HT+NdqOx43S1wjbJCUGr65IoROepHnSh7eh6LDDemgPjhsdyTmMOxchQA1Ll8FPh/5IU5hAm4944
+nOJ9FYUtLCGlA9gYrEVtXvdAN7+9FLkj9YNpzHYOXnLh0FJZ/UlIxObj+qt+IdbM2yVS9OL2juB
wEZkrgOe9PA/hSfjd7LbMflh8ok7kJmH+zn25K+mQ+PGOvS6nWqQjvOq8osWaOhSIGk3cHiCVlLM
CjG885vZ3MdxhuFkKHckIpBI96jyJM7e+Z7a1+5TgmCtvMtrZoHdBCW2H+mqWxM2EHxjOQuCEdl6
+MdmZzt5qlrujYdb81kJPNBthIpsQWQ/NS2w8C07usMYJQarvp4Bm15dLXRR+64zuJUlfbEa5eKc
4mDtnSVvpsnE40L0etzrQmdl8Rc6/smfOPbTifcODw+mnw+RmE2z4+H1j+qCWXPQBNqilVZwZ8pK
Urxqxs3+mIdIHC6RG6vuRmED+amrVCewW1+/lMkycJVAGwcxwkvGvQhKcRCHIAV0scNfmZhTSrZZ
v4IKMFWSq4oj0dVFa8SwDW2AFkLuGtQdHhE3Udz6ZPcme1dirmBhTAajAfXcTDTaVhwgi0xbALmd
e/KCVAxtLdLHr6+vkmk+0t2dVY8lHjhgDSb9nlSR/xEdN3TOZ+0vwv1DP61Tt+PvYFqEExK1mBst
30/fQtJyxN4dFlFNUBcOHK6mbBsTyH8k9sQgf9JnUDyqMpzdehkW38JsU+tZzVA4Lh5wwh7EcggA
vzKYcU/1piHIa353NleVqDIXyK3K0WN8Z0boIbnu65r/orxAgvej+lshoU/86wDT0cgExoh4a1Bj
OFzJCH61S6LazHelvjEw/uPfl4nqkf4MfZNo3T6BxZG/V4gC+j9tF/ns2xktq+GsIMpBpeNopj5v
dXX0OChudqInkeHjopGKOqXC6Zrl4xQs6vQ8KHaobsX7eYd0lykSBto+TDxyUV7VR3QNYoNbDxVO
ucCb02lHyZAS1LoOvI4gTXKMVqXyuJOMg0DCv7DTh0HQSUuyUZqP2j0BueymVcBRpV2Et2Xe/2TW
2IJyKHVH2bHw8mwo3Nio88GTtrRuTt8wGkcxdk0DvyhZ6kpzvUQDPMHdY64/WFatYGU0iyMqWAob
1exIMCxP7e72vf6DqPM5TV3fEwVJQ6rfLV2/jS844R+Gfde823dAwzuyhUjHCs8K/PqknSOCQoYG
qeBnxstQIZco0Btp48qBJzWca/OlKb5L0EIGkYMQ332Yw/SSwVO7NorjvflFX62GpByztZjVzC91
q20mVxIVAZKeIGMrIwCJCdAy7RG3qRugp1eNsDIllE3azgDXaMi0K5PtYu10m3FxZ5K/XwvLeqNr
AIKsYVCylYXIQWJXVaA5hq5lu+sSHdbIMuv6iIrZ5PhV5MSIU5z2jvhTLcDVR+zzKVa/4vDPE8X1
5LKPDCB+8oWzS7ngD5wK4/T10HTAlj40KSKYJXN5aJjwwLN9CtV2NhUn2UZYju7Yankyg38rb70E
1kA4QHNaphjlc4EP3MXX/7JkBXHCk1d4Y7RcDE77l+w5lbH4mtP38Omhck/OIe//lRU7S6vp4KVr
d9YxMIklFHuSvTJDCuG0V2iVJbjJe3KbLQZIeD/oD5QaPOWyw5wec0yOlO18rWPhdnUQn/EFKRJm
eHdoSDrCoSsShPg5jddzCqd1jmDUpeGtXuIZha0JWva32MB2qx4OH+oRm4Qgl6h15kHhRiJpAra9
PIPv7tg9aW9R7LLY/yQOG9jWvrS2tx/YmW0ior0QTHnG/c+d+kKkZppXpjvet3CkS7J1TTQ1+cIW
QoC3Br1b6oKtytWy3mZpxk9FcQmufVaU+e3viebbGh3v4rjSIPK4PB1+hdHxwSlpmAhq3RwS7C4N
nhUALP3+B65hbO0OD7y7W9RdESULu9M2EMyIdwAiWFgM5y4x0qIVGQKpvzQSp+cxum+5ZvJzz/oi
ZpTKOv92t7NYufQ2QzrQX63+p58hvo5zAAzupU9WaFWHU5gO/ua1gRdstDNDzVyWlH+vAO+N+S0N
G62xIyYqHlMelhDG75+UnhgywWTUG026/8a1Akq9eCVDd8i0/cjxC058VDyt0L0KoXyAuuvy7nws
uwTabnI/3Mpa6aO5EAeURqTKDhPqvW0KyhyOpasTjPwAwDaRkryv9ss1BKKbUgJ6n8ROiEOPGY6w
eokZ8AfGKzMaVSIciFM9jOm2qKKtUYHc63o3oFQ5oLJV3cALD1wZE8kl2dktZxzIainqh900+Q0p
ssrW+ElBgkGB4EkNmBQJnANzS/8gKoyGAXoY7mllvj9bxkIwkl5y25K4TKM56YW15bHfiTwSOVdF
f2JBjIGAvewaDplF3Stn9+e1xQgmX3zG1B8XrIXRwWVZgLhGObzPUnFJ6O8YUuDFNwIjlflW7v/i
cWQy/Juq6ImCJpWrCIqllFd0lBvpKLee9dkK2gBghCi1+hfWHUJy9ii2EX0DtymLcMW3VD1Pq5Mw
mHYRZTtY9OfFyZjdj+kVVRifldEjenqVGvXu+e1IxO8Ib6vgA7ptW3p75nFeY+B2yr6TaCbtOVwN
bVbvLboMpDO8wVzdfhCH8szcDT8ct6t9a5XhlQU0GvEf87THdRpjxQFr4dvTFUtb4MUK4ohV1xyh
OqEAGM76ucVHZ6il9zoXF0SILy7xL3Se4JxfGAofEesWLKfg0bttCm2nBRXjnoCmoXvM4kt/Hbgr
BaCAvMOuqiVfxcnNfYo6IQsBfKx+PTAtqywwukKKTBJw7E5crO2y29gRH+FIqi9NNglNyWmb7bsO
5nwQCHCYB7Om6My0NZ0B5EZkYROg85mxoFCvl03IHrFkbXqpJdZriwPWY+BlyhCyBCWdKnsWOasj
E2ZGB59ZSg02ha4vKL+lxT9eW3QfA+bF5x0PaiTy5OP8RohAxhDYYLl3i77yY/Eudyz8VzTa+RQK
f2HyQa5fd1jBOBujteZSiUo/+6YNssZGmj8WHj72V6aDnh3ChjHqzU5cmZzLx88JOOK0eKtlQolM
iJOyIy+rq5bXp9q3x6GbOHqJ6Q+7bWHCwqBPUZPEK++NTS3PxqYp4eF/KuILGQaF9Wa+KNP0cGQ1
y4uLl6cuB07NGqyHCXcIB3ctcMGXon6Ust882zyob/520nWZ/ctCnCIJ1skkjaX8mrlNQ9TNL7Zb
i8Kj4zMZMIJzQTag0O9l7W3x9tQyPMWXwsZRb+KTxNCmp7VNNQbFHgusRyg1dZWj5aEcJyYDPs0/
L/BkKmHIg3sHHPemRqKWvNvVHY0dSjfoB2NrEptKPmjhIqYx8o2qsLrAb3oo+riHO8u+CtHPX+B4
W8eYstz4Aeu6gHUHW+zzoB3D75O6hllDeVU4egd1n6yZ5rC/0Kyd0aEFjog5W7OwuuatQR8ICqSN
yCaMxNxdBwjwYXODXT+rnJ1WVV7l1uzaRFCJHVGjFfoXkscnLmh6DrvMTh9cvUUhTd2YRHMVo5cE
HbFegt+ZqgTS6fSyd4yOnW3sQ5rnn1qGuajpPrEjQ0oIgQcU4rN0BvMUY0XLRvrr+tG4SOdVIhSR
QebkumFKR0hpdMaqWuM3X/Sl0vgqZE2qtW+MN3deBDHW2P9V7M0w0pqtG7OYj6DKmo4ATlHWfFH8
Yb8lcynnlrelc8j95nEufoC03nEVyE9c/BUZbY+C6/SDiqKrglubx1Z6QTfXjJK14ZpHSSLwvGof
Pk+HiEsPhWEH4jVWtZGRELL0XYbmhf/df2AjE1BpJPLRZ2sC2+jcZxpEpLw34+Jg0yjU2RinCybi
sHnjs6ER0cRrZUIeZlwTEa70SYA0C2f+IUgTQBHhyqKgB8jx6HfxPT5zt6ySsv/64tRN34wGHeRT
HfMp+rCsRWg0P1ulE8jj7iughmQRaiDTfCPVRU65Wghu45ZIY0szofq35oIRC+istdOWQVNePwGq
VNOxsqxIcSHz2fs/QBT7+pNk6Z+h7Kah7CodeO1u/BX3/LnP3XIQQBR5anNUY8mSnP1AYCPNn5xp
AZwKaB+vpoxCf5UeVUdA0ZlDWx0hYHNsnEGnV27JYTw4hVebCRkK48oX4yZfyaZlFb6/2lFVRpRD
wWDtW5VvIlGYv62nMkBJR/tpeq4CMV/KNbyk+Oh2/Z4z0JdUUYwwi15sALbKg/jELvV/IYaZ/bs6
pxvIHkbtIYG7M4isEEV0rSzS8gc7VPLQfRiDCu/RUbtzfkgk8bsKy/KhEB3b73n3XcJ3x96xpXot
uD2VmVhxidXTLSAws52Gstb6rpQPNV3f08Bl7JgRCcQTwtDR1oKWgFoXhsbNrcLmwE+jxqmJfmtA
wbPLVG5VVuZOxZl1K5Qa/MmFrJz7a/PNCzdZsNKpr4tM9IliAGOqk3jYcQUww1bYXeH/67LUVytt
bIAZUhw7KReP32gfBg3rlcJUC+Vv85LIoGFs9/3e3+ZXXKObx0+nLdwuUwrNZOYi60/s1BiANspq
6N4XQpL0bLkxpfpSwAjwDztpBPsa97L8c/Jrlql0lggkeizq01LUmbFPCrpqUxb+UUFO9mLHxJXh
ZQ32W2TBi2QCbKjnRkuMsZtWVGN9JPl0Mw3RHAYLsQkQGIa7mzyaqlpp8691+st3qsuIZ+cgLVse
QpVGSQiRyd4ODP6GEfKlgN2ru6JFB2whSf/IO9rcWkKhPoQjH1VImIXR2rtQVXeSt8mHsQYIIeQM
/H1+a7mLe2ZlnGDENichWhtwq2N2e0x+iW5ehviuaEgWpkA5y1TdFqnIU6B9knd9sJIJ/5o5pV7j
Y1sPM5rbvfv1LAy7Te+BaZCYbQGunRSx/2gsFrdYA6o3gXgUlBDvlYyFwnfS3vEgX8v29g3PlqP4
yodnZJ42hGqjDkVrVfWvlpmuzslAXbx1OTFJc4dRz4kya+85qCEWc6kMYjEIY3D8GD2WXnfzBFGl
NbVfC54cJ1CR9iJfBq5kpdF7gix3vRConSXcS7ppga8MPsvOCu0XdAFtBZT5XhDxZ94sj7d2Dvg8
S7Z9xqz60lDfa8PXgJ+maE9Yb1A3KXBVKVW5k7MSZwxwDgle5uZF6D3+DuWLKGEWDsZRks6msDbh
gMDd2H60So16VfupufsPQ9iQv9ksnzIdv/eAQiGS/HRISJAFte4kEslPzptVqgwLatkNVw7M+y6r
aWuS2JDJdadL4F54yh2j9OQEQtk0XzNeJDTxAhvkeRk00DpYE6zFDz9SSMw5R2mjk1tljIrIcFkl
NoPT4FL3kdZPeny2YT67Thzs9PmXd2v2SlIoOuYgdDaZ0aL3JW6mzk5PJHDzIzKE7Fbk/YJPLm7j
kB/wbObN3JLs5+rpdP06fLtBQsF+K3K4tfwNX1RNQuE/T1RctO+pTh/EqsM/tKQz31cc8+3qt5SR
ZlxQynpZkdH42gHvigiHycD2+w9Spa4joUXWES9WrkLqhnNcXqt7cWWc8vkGiB9FEdyp67nqpjyL
icWizKS3Tdv2tx4bPToVJI2baF/cp0af+R0K1hJfJRIAjLXSxrPDRrAhhtvrd+EOSUAHDZf18DD5
o3W6njn/jkQnoy64LPS+PziSrVE0h13woRXFBFoi9ZhuYozsbvRpGpDc5ZLVV2jvA1aipPdfHRVg
Fy7WUEWaoO29MQwUoXj4iteekoS9IE8WDbC7+Y0dc8FItHOr/k+FEbA1d7vBNjoAl/ZijUDG0VES
zVYPsoPXyNiG9K+kSMZ9E4LilYDSyE3C3MK4ilCcWoYhUSIsUeNA3YdlYrttRx9C3T5hy4ZQQcCz
jrAhLPLONi+qKkAMi29V29QwFKfq54GhMuQ2k6bYDXZmPnmPwfXztRhiCyVuc8y2ktjG9vJuYbjA
2ftnvg+S2YxSd3HyERC6QFrQn8ZzJF3QQQaRnuIH+BTyN4U3qKvMDHzg8OjCMpE7d1PiIiLLYxgL
SNMGJpls011xEYA2SS9A95eR6UBeHdb26Wz/n7PNsv2wHT+X8iyQMm+iuQqArGLqNtx/oYyq4OSi
q5ksWyuGvoZMg/wCuTJaYjBn0YiTfeRE+htuSL+04VD07aU+y3APlbEPUFjN0NEja4Oygv87SzSr
ZK0tHwRtGLmQ5LcuwPJSocaO2IZ8tMQwkAttHxdpXnJ8UuzHCIYgpaHvduslxuSuVsK3WYhYxXCq
ZedqzHxzcouiF4JcWxfmRSCUhdZpL1cry9NFzqn4/jM94VTfukeL7slnabri9eGOUDPn5zojBNjV
yhM2XiafEY+/aIYOCRZ15hT89FV1bZnSKfQKFOaM5Q4XtdcRyod5Sc3UBLTugCgJVvcrTOS4Dk0O
y1zOeixhgouhY6usbbvJkA9SEReE45f6eCPOwSvcZAnBpWTNqHgFmUiz4ZtmwGCoUrZsDwLG8Kf3
mUAZszgFSFdd9vHNQVszeHKhscllNa8ht9KJP/Yo2nKQofjm0RLs6baa27P3PN0pyVGnRuCeya2I
EFOvx2ZInWLMiprBmFOn8ftzkINPtfCwkS39t0eQRf7mfKrWuy+JCKWl+Zgk3D4G8LJ+jjvdFEwn
24odw8npj/6VhmC37mTsEUo/iMfKhsQz0VyMqBLi0e/9bZ5pIBbd6fn/Cq9haZFsh45ib54X+VBc
UIt7tcEGnuX3RJMqqPUfHAagyowpasMdT3T8xsuHxKDo485NPBpycfm2jLRRHphTAU9zDSI0bPVE
bakdhpU1UGXMX6M/D6IOKrM/eduDnX2eMzEqXqlpwhMaOB8Ie/9ZICSRLp/91vbACiLNT2z2kIiC
5G5M8k8doTXVU2ske7WteTOADtP/zryf6NJFtP7EoBxey+z9fHv48TqJ5JpMbk2LIwcU+mZGeFdh
c0ERngx9Gtb6tHniX/J94tNzznKXGscv4x6lGFJf1ZTAxmHnP5Zndvw/NaGa1G+n3dQrNYS+Au4J
ItBb0SRqDTNrswWGfDmUXrdG+PcmGUaYNxgcjPKGwH1o2AsnNzw08sEOW98mvJeOMlMjPSK0VsCd
CNMKnmpMX0gXJ/ey4dlwRqxFK7xIcTbv/+jbRzx56YyYTt3SLs6KYhS0DkaSuNpUAeMCRiSbyiWE
he9k9lm8zDOQzTRqa3oTVi1kfDF5jnPmL/1DujK7wti4SIVsTRXkoBqc98WjawlsHoWt3OAiYL0a
lDlYqi2FBwViwGApWVF4EUsEPBdF/omzQrCeSQY3qIVkp2+pnwNYh6Dw9HO0U6Di/SC0/stsBkjd
u7Hhhj6FvBV4XnXySlK+MGMTXzYvuo41yOh7wykMP4GhrZekkN3hzNY4Tg4inGKW3mT1piQI669V
J2po6qEA1N2mm39+5UVlrkCBfuCsYWzvHpmdDWB083/kOuauYwihzd+RzVK5q6+aKAoDDvNPo+Ev
Pa/zvUSCOfJe+wm0tKCeyVnR1/KX9v03KInMRj7nAeHFtjCXtysAfZoys6B9W6YxhF+CdR+ouqII
dgyw/RSenqqRfiqZTrTKKUGk2f1zEIr+iB6i79e9tjt+qYz0AWdHtnQfFDA7Fkkc2x3JQnWi5cJj
RXJweRVLSxS4x+LfJaEhrFkGxECbetnw4f9UZgpV7UFIjcGZFy2fX8VsG1IULam0BeRA1mc3Syuq
IwxvCz0XHRQEgV6rVovvDvLxTlNhDCnsSwgOrdrNm0ZY0e6DkyXiEMMy8ZotJgxLgUAs40E6+hrx
gDiwuHUFCUv3NvDyHZK55Wv72ULUHNjusFfmO4dbRZEgoKOuurSQfhoSvd/5+J4HTG9ymCOT9/nG
Jsyn2/7/hEUnvoFS99hpccB19B5Nfgp8N9RKefKOZ85gv6uyWstpek3UJt/6qVu1pqQBhLnz+SQ4
mHKAEolXA/rvmGGO+otHgEwsGlIOjJf9E7sXJtg5zU7f5wCr89OLs5bHrEMR426fNYn/2EUzV6uX
uA471nhsw1iGDWXQCn2tRoJlRkJSLFZVpeaOs5llUyANNRhO+H6Qqy+VzbCgcKIuoNfHYQK4fqZc
kb75Clg2nU6WKoJoCd0/r+TUSKTIxVaPDkCJJ1LAGSp99TSNqLbZ3DICM3oKQ0rQkhxbl+2giGC5
Vkfg1QdzugEnwbJLR2/VY43zyD8jox2UUaQTAGXfIgKPACWt5bacrO6BhPw1dJ+pN+3rT4zfdlYh
VthE72ibiWrUyMAOBzWioJW+Kr5ruLcrhnPWYn3CkXdsjo+TyYPgIr1iFJ1/avpEdWEMaTG/cVLA
tMHyGuK/BnBHF8zIWp5SG+pPmeHY/DvW7pShfIljCHiQDkLdbtvKLaEbTfxJe7VVakQH3i4UIVBv
r219JsHlka+A/ThqpxdXbUB0VQyJ0cicxklHwlymZNBTymJSYIDIMjKt9dkt0hP1hxIH2adpy4GD
I36zZ7JhwqT0UBXKczjmk26j8kyUKwgLGf6WUF+YQatB8tG3owIyao4PCP6bS/o/kkMwFaYyVuEX
dD4jnajilCZU+TVJzzLvuDVyYh7MwncAGm8hgYwP7B6wdElI74b97BmiKIE/r/CnsuTD3H3q7wl2
Dko+kVG9WgqQ/L2DV0GGuh/VAM7D9BlBBxRg6PVq+UxbPwCXF/l9sFJYMtjbtRBj3hQEGJkUl2KF
cUE69crg2WDSYv2XnjN5alKrqVQpHVV+pY3eJFf1RPq/XQmgtpNw8ctxfxwxNESaGd7JnSKFmlly
zZSLc361IZPu7eHJt7f4aJ5TYpk7cteEYEkPiguWDgMnT7eV6wACXfuo6DNcXiF+DxpMDyM3jhq3
zfcvFQ/WNi8ZIx3qFM4TrXmqWvPB2s7KXeygDJ3L/I1asbl/Vwdk22FhVZU8dIBY7af6M/57cWlJ
5D5xVQJyEI1q2wO0Ua4u/2ViRNjvwyoZjMKT/ZpWhiM7+TVny+JKhW2jSNO/b78NsL/rFzxx98M1
Fvlxk/ePhbLzej/FBxx6Lp2RjEJ/pyG5Kq8f1fYBjk6bIDfpHC7RA/5ewKbtg3zK1u/ntOTI/m+C
XR31vyXne3vz3Tw/8LmZyBz62NJc+A1ZUdq5zVpWA+LExTBC0EMxOh0ZWKJNDFCcTn20lR/44uBh
3GDdG64qmNdViJZ01QkBdB/a2xsyL9qDtRrmwqfG0w67+608dCYMfgB2yVFhcn8fsHQCycZCPKTq
LDvGXe1I1aHzqFkAbgWIkJ51hOZLhtEYvXc1twSUjIkQ7Nk622a3Cr8nVSSr5UY9FWgW3lArVaPA
l0egE4wado8dSI4ZPt5sPNY4faQbag0UyloYCqOLzeGfVsOu9ucIcdqnXstgcfl1gD2LIVa009uq
fbK3v6jMKHX+G9RhgesPzH6IZOs6vgtqH/KjpYhW7QqCt2EvEkQgm03IbFc2Svy2VwGUA/ngoTF8
n85h3EVLOp+TLyxgyKqJmf+zZWCyh1tVd9cOw4x3Jm+ARendGhVqknSPKnLWc5moSkRfAdqnM5nc
pB0KzOr52GUT8zJzRcBa3huYZvsC0tuab3fSyDs7ETyCMSkT0de64JQj5OT/bU1//zMOe2qXQIXg
QWvycvPvAvJwzS146AiMQBv4EfQz/wlHBziQYLiiB33qZ2c6yy9IaV9Gabw0F8KNDSO0g5RD/Q78
UjkdD6yQMQecCMhUBdo0xwjOq9y9VziguFxHMXHhsR7VhkNVRxqB8UI/p78BdEEv++0P9wIQh5NI
20u5MMEd7V9XR9DmJgFTuMRhagnRNIPgl48aj3cau0Rfe/2dqvFy6QLHWEFqnoMvFh+ZzPbd0KEA
FsMsoOqkxdv3bJCtKqjtSoTFz2A8muYVh2MmjbYyxVeJdWN50NCW5A2pMwXtTics/0J3NhKagqIr
EBByV0n4lPhoKFCDn1ECgaD+MXVAYwo4QcbSzRiksrgAllDrjBuUp1osy8VmxYNqaxCL3GedGqhj
LbTrr/GtTYt5qxgVKlulrccCcSgTrj67kH/1TqT8qQncm39QZ8xzUhCESJ6Z4po04T8x3q4cv65e
XU1z0XYnDH473BItY2RTJTWuvOrP153uMoNHQ7+h/vx8VLC+a/SEv8/B/tnboobSaw4xX2VTPs4H
eBGcp1+QAKKXk6jh2hrdMrsGNbiDD+x2DmIe4XG4wZiBOsMfYviz/Ib/0RsREJ8koXA1ZkYgARuw
q7in/m+CY2UwxsznqGzHu6uC3h6alKxrKWcnGjPEJtLKXyestkJTofKpe6OQyMt75tQutTgrMlLa
MZK6XjM9cOEYy8R1iRl77ZCY951sPUFMi5AHNYBPoEc11b3uMx1OPY+rA3zP7hOTxmIEO+0dg92J
S73VuHLcswyu/uAmt84l8DJJ63jhMiBUPZDVyKbRPJtNvad9dD5ZdZYctakRhQQv7B/9aLPxzjuR
5iziy1VVV2+koJKAQFlo1ypPe57uHBIg9xVeb0zlfYzxPnXyXGYRXATeyHZ/zkdPsFVwIlIybMc/
cGVqnk0Shded5EeTZ8GHiJep0MnO0FgX09C2qgDTtCgonMWqJF6Mb8faoaLZQT5DLiyCct9ESbJO
brwwSVXgSatmQo3oGMJ416IONkb0nh8kH76Egf9yJBbJsXnWBkaEPyFLAAA4byA/MqLxY5GjflmV
i054Z+4s2IUoWkPTU0qYGusHlYv+9pxDM+fHdUgB18B3bJsT9NKJWel+stivqvt3M2iRp/I+pA3x
THSUUB5YXilCCA8IHcrICd4U3rMqSMUTWllufjRkp8NQy6on378amfGizetKHoR/5V16KQmIErFI
isuLNojnoX4StwgE+QdxP9l6oWJ2yDkrWRwdWKF5EVM9S82FrT2vjrFgzlhMWRKONSNQ3kwbUEpm
OJXdL35n+2DbPHGP3CQn63gTdX1zpr82KJ/0FQ1og/o1noJRhQZaMIXaKvOFcliqNED7frzGS82+
EWpVv95n/jGcbuRrErf21MTfpvjfdl2oxsFuvK9KA2fW0WUPBQxqBsLeuo8cg6QiZlaOlKIFlzWt
TpYOHQ3eTd9Tny/wLu4Lrg4hfQ1K8jGFcXg6QgtF9eo9uoK3QVylDPxYTKJPcCXvRvkN0hcshota
z7JdI5Olz5T9SLcXm2v1C/R7mnvRaIrCxufJAVJYqxnncUpNHEfK+TnaeHWfVC4mT+Qy/Tufr8fK
VtQ7n3S5/0fU8fHKDBevHOYw+7EWodfpahRmZIAvYzF5X7DUG008CcBWmGfIP3pAYjHuUBzzGma8
6ozPzxrto120zDJNtaJr+kxc47ezWFlq+rmIKI5tr1Bv9hXCTiiz/PuYOJ4TZBgIAf47aQ0QjBfB
GBNWZKPjQIHzFQsTrfBnpj1bJNHjaOYZxDHMxwCJLP0V2yI+LyXPK8+Jy7DA5sD4U4vfaZGMpkDZ
Vb1ErXhGySCPk5lYIksQBS9XlQHi6y2aLinR+5f66IMDZL1EIUr4S0+uTtucF1Hogm3QGkG/HGcT
8tVfIKMZ0+V9o5si/dR0xrf+XXIyqhIF4h/qq0lSpFDT78XnZ7s7vuySMOboxOBu8EteFikjjncP
mQCgquP2uDHNeI/nGcKLvpq69yX7aD5azHk2widqfeGbaLGqRopLD3vo+pTtWLUwlz22XHHmkEfQ
svcfxgvl6El6S8AhTCri4lMep35gyiTHyzhG4MIzcOVhc8uuHETszTqYVEned8GXIhlFK3BhGhOa
3U3owHfV5sT8BXgcW40U+535PPnmowMKrnp0Wdf+S1rB9Yxf0dCRQCmfEO3LaLLnWEnkFIH4PPu8
qIiLmJnEGuf8YoH31c8/YnWZDHou5QVeJTgpvdDo0ErTc6MzrvGUQHGftfB1RyBoDwIrYsGvDnsM
4cavcfo9gR934TuBu7Q+U+bItE6u8yyAl+xJ+YllIEtbNOBwC8movUGZh7woNPXH4OZCuHNQ1Ohd
eo6cnn/k1yffBXfIkYjtdwXCzKZIpSu7OyxC5GZpBHyQ4fWrf2pgJAc9DEWqOX9FNbSZoabfI2MH
92NqdzsYsxCJBG7ng2OcmbY1Hov1d5Ke+4bV4kF7nwwsd6alvATLvtPxynLZ+aGArTtcTQpqNh2M
SN5/ascM+YP4hMjs+MqCAix2SNcFobUSlQ586VUDIgCS9POcCRMwl4I83uwJsx2fd+vh/ChhNPAD
3K4ofKMUzlvcT9mTuIscv7fKcft8SzoGH0uUebDNWfGnJi/cL0ts8yGllhnYKV17pVqS1JN1ntws
C90meAbHKiWfoFiO0Slj0pR9ewNryFC+/YxhbEjdLjsyE6zmk77A/p91dMHcjnT2FLBZe4bMY/U+
Ak/2OnkQewCGlC5jGfTy8EICO+YBEAXb/HoF5QJHeVpVw2l69DzPZeWuWn6Y374Ghp4OL1mtcJbf
BRTxeuScGJv9V6oi5Cvcpn9KKqlkpu3OLSi5qAUzc6NoGELH2W8XaHA0qNqNwVWnbELKmuELZLz+
RnQmTwpQ96SrpunjZgCiIf2FFSt/s/i+MESEM69+Weio+7oGV0Sw6cPNRjr/WbVqSCxRv4S9LTIA
pZZmg0A3wHoCuOAjfCS0VgIUvRrxxinTPobO9vaM1I0SfnGOyYfk4nKbj3RUDZjgsVYm16rXHPDE
kJmGkd/YmxXhgC11RY7KDah8o2Tg86kSKbVzFyI7ivyWHgvkaGIagFJQO/bwjihT4JhNCwntrENM
ci7Ekri4DXCewgp5+TB9MN665I7xn4wAzZtBgdM+XznGTMS1u70CvnOXL8C+03pQUmr8Mi6gq3xe
41aAdRgOsY+P/RhcBcuDkWwNHjABvig/UlQ0vWbZ/qvncINPuB8L0SK9v/EYkb3IPxfxCJODvyw0
ybba2tFvI9V8GMHkO4XjO+kKj9ewt2sRtUvsSspnPECRLck1+y2xclM8YZnywbZn6rpJX21odB7e
hXstPHeEtM5OYpwvTypnFoHm1L6Ih+WN3RbdMSRQlPFd1u30f6OeSpuk+tXKEZb3tW0t4gF03vca
gamSiaWjT8EFLDtbP+p7xh/4Eho3Pxhv8/wdtRKE3/H5zzACgM3ebidJ3xRQ7Ncb2PQlJodASB9S
mqvKAE/gJ8XNTQl885zQCwiBIs/VZiO5l53/Xys7GIijv+qPIoeIYv3BfXS7FPQ85BrAyKEjn4md
9s4xisF8n8S5ne1AaNOtzVcFtY3wtURLOhtx+dmxILwY3mpBmreFwrb3ktToH/M9RWwFY0FxrP85
/V9yCBDg0iDTZkLDv6kGyqFzRH2/3KeGjA3jcV03t7I98R1R5g+3hfIp6kS7xys3yrgtDpnQu83u
rOiiT5T5qQ/w5IhKNRCNVP5ydbdoTj328yY6PQB/1sabFZSsSYj6EwTExtEVp5zBSzuAL7RzuCGR
04lH2CoLR9w6VRPHc85U9JROIJtok/P2bo2CTfMCs8i1Lk83nC7O6u5aKIJheUWafbsqWYyQxKXK
MZQcH+CKuv/oXKYh25mPQwdUtEt+ItJ/i1iFALO51Xw7mtu+kXKwG2NdQMUsAjvYCOYL+w+gHyAc
sop0DXLlCsdM3PgqEnFvgyQtEYToNGu7IbDWzALXZ+pxZ0Z/v893PFjs6Ig+dldAMTWBy6TLRtsX
rjqCdsBcYe6KdRlFJO/WRVIiurhuBaPcbJt2kpga+umQy/UM2cw5houiZ6rQge9qXZV4d//9OieE
yAQIMPxB9Ip28K7aDYVcDMDq1f9kfGtXcAvwXTmO4qvMvHVF7gRYGCnhh1FDVcXCuO0GTyrLUtsK
TYcIvr4oxlnrrz3tq4RuA9UBiuoQmZK91VDkGdpKLtUB1pg8+rsZNsuD1ckgyH/LQBsiII70vutB
JTsUoVt6eiMWr8L3mZ266TYr3T2tA2Q4PSfyy9pJNciO/O7PukOE/SB1WniLsFCuP01yRbCVJbrI
QWOjuY8WSv34I4Z2dcPb71OW+2wAVL0d9gqYYpSi3f5MhgRx+t5wVyzsLOERKWmTsJrXQnLVTXyC
uLcITLlb8ivjIEP08X0UnNQ2OO7Xs58pBh5qa9IyyS4/sSPIpRr1kA1YsripKW9kOXLCoafrd/6T
2Jy7Vu/R6k8ln6ooIDtcAXrOXz9eig/vbNWj8KnYV+LnD+VqwFUt7omzEEYIa/m8Sv5kVUO8Bo6Y
pCUKkG6N36UYLjpOXmmYOGczJZBdjZlav6JW7lBspJPrDmZHOBlt94pcGHEVR85ykw1vlRB938Od
2rlkaQ4dR2Rjg36ZfEhr4PdtprEvIj68oQF0XYOFLSqAjraJgNjMwJWL0rZw8h1aWz586t8zqgND
0R0ihnkzFZQM8bac0sBD/Ab4YF10B3i63cgPwDNplYa2vbFubkKctjHOh83wiPqP4GZFpNUaIElk
swU7HS8M1eltaSIXLix6jxfQ8770/70LuzKn5wba4BtvTC1Xg8juAN2AK17+zgXGBANs2mEeTw3k
nFjtDZKwajfygUKcGF2qmI+++BrSbabOwIUcchdvOOim0gQDC2RM/pGje3qcfZIvvzN9M58leayn
EmopR3xEEWo+TVX9ojKT5qSIXK0kJI57LNpNb+gumosNKnOrHXK1tpWREMCEIGjEyanLcw7JD9Nt
djjfqLHbFhScih4O054+Zu7lFssEcNllBHaU9TwLYQgY0AzgdY73TdwvxwKNXiBcYwVJSBmilp5H
nSsMxO347o40R3jsLPVNnbo9U7gjXhh65wqmH3LopJuiUif5k1Hn4wmeoXGIhrLxAUAXkLJT8mZs
Sd5ky0oxNtWKUxevxe5uCjzgI2OEVGoylBN8tJKV377pZpK11kuV9PrDWlSRy3gxRBAeO59xgoMI
GY34M5qOgbZZrOjX3hZMVFKArTT1L/qFhZmdaRFGDklVh4+xEF2OfqwrA0hxGts6IjuS9unzFihE
Cb2g3fmkXxxBp6c8vOIuPDfzHaHWf1PhWzI20WJe6B7Yba++75l1HZz4oz7/gm9nvR7LMyy1eXgP
e9SL4QgO8OjXd1VVx7g7nTU+QJ+DhZG6ON7msLcuORikzMfYvSFE89J8HJDQhfywQTThBW6yu8Hk
iUQH35T6F813kS58haPnaUN5ROIbz6+45ylHH5VdbF/QKBTfpXHhyMV4SoBplPPMhhsKlYtEKIX6
TRUXAhESgKnKXjiegaMgmmrE0iE47VPB5PhyBuKv4p7HG6smcit0cjj+kyJerG44JgP5qshaPFip
8G2IlD9o/gZHuk3gHQBe1IoAa9w+qqT8qj4hlBtvHbm17DEBPxUq6XvmLdzXPMceuwjrRqtH56uS
TRX2URRdq1mModaJPLQBxNFNq/UGfs56Kc+CoolXlifyjYbAmZdKopsdBhzldIfs0S4+hTGY4B9X
aPvd2Nut3b7MQmIlxCP2Qj0kqbqDl53Elc4iMeGN6Yu4kZJGnFIXTvDrKSqYFin63VxAQtwC/LW0
knZt+fRqrn4Cx+V8K/3nRQeuujFUKhrwS3x6ajxW7gDaJazpf8aD8vvmYS412HAPKBUV+33H6CJw
kROllBzpd2wgNzHIGcPJM7/TZZdEcxVCp/UqkupZHJ/IV2B0YYHXAPgv3RQikTF14X6h03B0JhSW
7LO53WLApcH5XfUvI01QjgOT9wBZFGcZQrNQs6DCxZ68R0QoIC7dkG1CHCRjTW8x05P15JB8Wbip
lnJh/AaMt06kr3EMg+1rNRW+DHYs24gcXYVyLTfbqVAClUw4LBiY3vpwaWQheOkfuNDHky5Ur6zf
zuKT6KF+yE8QwIBxifqR0mAyCQeHiKQqqPFhYzNMAozCukJnDKp4kTe04wc2vW85zJe+2bnhZCLI
v1pmB+LGLvcIdkIii1+G/ukjzWUS4DVQ9JQz0c7dw0Ru88wQE3QunEOZi4SwH35CS13JxV5xdhZM
4ZptA+HD1n7JE9otFw6840v87a24NY+sjSClDnNC3zXNdW0OTK4r7e8BghK51Qyz21Kl5LZm8JmB
bwYu2cSQbDJlvHmE9KJo35jMxonCmpLEbHhDJJq+eX9M6Cif4bRJGoSoDBT2q40ozC+tT8v897DK
rN3AMAmfgi4H5NzzSd7iOkfPaJnB/kxfsO3gdiIbaR6KdsEYKCiSx3rOkKb7AQLQtPs8tAejR379
BAMFfXmV0J6EFk2edN75GQ8ZPqvmXWgi0W90ODQr96AJE74ZgO0qc9o10lZzLc5OcBZmhU3hIZ+s
TLur0LlYa6sBoOEjb151ZTt1c1Q9pIYCvOr71SfYjm3+2RoGnlT4F+jEBkifsn9e0yCZqP06Jyp0
b8dzXQSuHl1ahtAPs0gGDjLWcpBYHhFa2g9b6qaeDhhqmickvlpj5DsO64hCRH811aUDrXfo60KS
LKzcUR3seg+debFDdOdS0TchRr31E0qGH/dKDIvlclw0YsyoEUTfSP4XCfQ3A2ssO8qfaxDaPFjv
x549z4V1FTfi4ZhWbCOIgMgUDUMTqxWf7uXucWa0uGCAEEAZycOag/QfcAq7Lk1jgi1bLS3cVhAm
ACMtKPm5LfZxsppjkwFO+aXbxCRZGwoCDEa1a2kwcZJJEIEeHWGN75Z350U8UvmIU8j/GsAvWliK
FsO8EpP94qyaBAuiXWKjsH9yqeLshx+d7hS0VC0nyBxK6qx+jbFjI10p71C/9CCtLVCLynfb9WbF
CyB+6wk4Ev9pxXFQV0+qo5UbVs38A22/2isyiapqZVzySJggkGaTZkBuoWImEqnnBpNXhTi48yze
ps/hV7UiZZSF4pwnJ+9q8JaKy6OwnKUET8JD1f60ArzgmwNA8FMkj3cdHcSTL+nE5ICaQOVGLqD4
WfSFTW1execNaTdvMggLEHOl8/T5MPO0dkP+6Bzd8FP1LqPXGyKIkUWKvVv82YXUR11NTob5n5bA
vULlG3Oyk6xQZ3gDoYHVkakChISzBv7sJ0/JqmfIW2Ee9LOOy5tWVSHD116YBkSbPKqswKrBJhHt
r4qpOcFERvBmYaFhOOFpO/fjoKtxJ3i5sDMAzvqDZ7VWcMnoY8c/kq4u/jF2TMsD/1l1thWzHyYa
LoyHJjWTygpugt9YADPXj+W96nZ5mAt8iUAGtGQMctYta5uutpMm8Nqlmw680YUFm4UyFhNj8RKB
9uNbEpa2gHed17odgaypqDqg3ukszBSXz3djgXpTWtItYsAxQ/2Dj/ZCmJPOmbAsvExZly0gWlfZ
gn/Nmb51lvdUXIgJRSek8YTlz36OZq8fQNddP2R+pnE/lLTXO4Vy5K0d5cSK5JxOTLi8oZvBnYjB
IJom3BZQL3kTKkbIzwLUnPHoXhcU1EYihJlVfE56h1AJCf+wduSI69SVTLitfl3yQ53pXxRfj4P1
dINO3oz7cFP7lg+5YRFQi8mcfw7BFgA+xQQn1U29kP+4DKY3DRUbdjZOmuBqwQi3f3Yw0zsYECNY
AgHUpUbR1Qq41JC4eJr5nRRYnucnC0IBZeGe3Si7TKF8BDvTvggwcax0ATKGoviE83flL7b2p3ss
6k39q8eR8LpcB1k1GvJ17XYPZ4dbJ9TfTNKzFfvbna3T0lJid0yLaFWBlSaSZemWkosuoN6hiFNh
hLx7tlXqLZnLVhU+dbw+mI2iNTEcv9AAOxpX3G89guFjkdpMDUszKu5ASzxcbZvJY8AfoMD/igY/
Mli9EUKPnt4vP1hNNBak9Y0QPxcLNiGYdynVQ7sKYBIKzuYBZeGuQ3wBTR/K53wHvAYyDfxl/Pau
U4eN9+8gtfKLNT18+LOGP7DhTUA9/U8bdtdGarmWkxMWnHeGk9sGHhNZK/20mZUJsg05e4ungxzP
kGxW/04Z/yIGuJR4kj2+rkMWp/hRQe+MDGYmnSokYBAJqCe8NmF0d5mXgsvo3pmO+wEkCnNUABKv
nAWyQKnk/Mbyiyjot2+eSKdoYn1cB7SbfBkG/u2/pknFk1D7STZH4xLs+SESgQmi/ayLH/+CreU6
DCDVw6DdvIdiPf7pIOXelHl4CyF3SueB3A6/XEzUfkckki71dCABsLfPN05c5zl+BjhaG9jgq4pu
Foii2OBPkzMIdnIFFWXmCMWOU868xb2uvCtlu3J+ou3IPo416czMlvLRfg6jouw/OKi5RiCs/vdr
IqGqFMJtGZjdqQxqHpiVoFFIW5BTvrUGjrFna13emVAScTwntnu4AS+MbncOiyq7biyzriP8l7QH
XKzG+UeYgAthpPmulupbzArgLYqhrbpfB81i2EK4iQt9UMdBf/U2PNVBBfkUtJgAc80/wYwxJI6c
Y1skkSoEonVIjdo3GmYc3aAUDirkoi88aLNL7yDt18UeDNjWEmpR3T0BsE2qoZ/P7w/LI39IrhOl
xwRM+jGQs33jtACQzknEYu2YnWM6iGkj7WJ1000ALaaTYZCzbg/evUUHtOq6MDIgno8M9ysIeGqo
haiiaf2ISQC74Nm+6RLXgH7rZNT2RlPG87Yw2n49/yS7QjHYAAO8LsfBNDmYDvAhGOffn6HKarPS
OyTX95o9Z2Cg4LPzIs+CCZjwUO0FKDe5EHfbBS9AtVL5J4pXbFaPtByGpPd4tM8vTqiG5oxB26kR
aBKWQC1bZPdjKosyQyTyUmqPBJ8V4NbyIANRaeU4HfVQuuyzzyxpy7awQkvF0YUGa0pvm2knnUe+
mBKZgYVACXzSFEwGBV42PL64MI8js/ds0oJDg86xRkuS0wTIa4x+hPAg864w2Xb66U46tJ0OicLw
Yz9uNqeNzNyUKw380Ulhu3ykJvaAKHR2GCq9oQdDx2YHrJ7vFOFYWJ45OhjrFSudtsEL50JPhtTd
nv6dM27kbSLdWnbLVmWZ2k8PT6S1qS8GbcZpxQfvY02fe9KtYU/WeVhqYwSIHjEypmnFQsAvhyLl
mr6T9doHCbk5NkGuDfDN1hTlBzyh8M1XwdWz1Po4uKS2vLCzMvfuWlJHi57jeh6ChRX1KjnKvVb2
oQDgJBylIzAr3VibsQZ47DjxjaGz+/gR72Eb7tYHSlEBgOjMfYXoIkbGw/IvJw69mo6hQJgJYvg2
hrEB7YrwBVOsx9sbUNpgDVBGWttQZW3XslmF8mva2QzRzXZRlQJXEzufI4TwIVhO3o0Sclz6f1E5
cm4jGYoBvV3cC0FWa0/76ZLDyqdJrsfi2d0Efv7tpcACTv23IkKdKqLoaJ3WQBf9l1ZdFgw/NX5Q
DSNANG/J3i9qZGiwu/VI0E88gRto6fNEL7l/XFRx6ntIDvEMRt00RMnkjVEEuoAiMpjOhdWOpPFU
VTTTZ0jLRU8hw4zT271A5R8ODEFvnBHgK7j0yBxOs2CwejquZgHMqFeI9KYpmWLdyPMAvd4uvQVF
Nc+VpAVMAv0zMXoZtOlniC0EaFPgJk+PZ0ipLypJEdLVT9nzSRpxvhiEABRyeepoEyEJ5s00b9+x
rX6uR+vCeCnUW4RckkX2fMweYSjhivXDoCyFlL1ib4QSB/E+4IQN3LE7d4H0K44xKsC+PFDYh5NT
XTq//SO+Qe0bw3/L/dj2iD9u9YjtevyFBxi58g5zDl1I2Nx16tUn9hEVTfb2llrzlm+pYsLfekfZ
B/QTTtId8CXEPtATYbHgVoNq8PC6bHtLwBYHwQo91e52ZsrZf86gh2VV3EVDgUPYgJBdPgH4qtvS
CZLROPsZvUDbT4PMv6AVmjn5ZUHSkhlecMf+GCThNYZ0/wC3/nR9+VcOVWB3jWJT5Cyp7oFKGIpf
y6EISYJhrywfJVgHx7m3j4Mcd/Cjb8+/saBG2NS7PYZET5sAtGd+LCEw+N7Q8oThldznATcH/AcT
joVPWZR4bAXHrx2HcE9yBbw4S+0GWrJXgmaEtLIFy/WNLrW6QE8q6ZYVzAJv0ddJhAvrb1AdhQN0
q7TkcCG1YWA1+GPd9nhyfIYWYRs8ykzp+iGMCRqKmSTWXtOtGIbEUlWKekhujWU9eMIMP6zApkxz
1QuNagmhsfoWEvwIRsHxbgVPqiNQrPAMaqJB4Yn4BfnSd6PQ4UYsAvCHgoVvJp6HCqR+3zxvPO6u
PG8ncd8oK7wEd3gabi+Ii0F2FckX6T9C4ndiyW+96EHXbFPQZjAbcKgyO5e7Cj/lwnmiI6IeD9Fu
pPAIU+JvEAvB0m0PoLf0v0GkAaXMkjg7zXrz//4cusbhzKvJgUzpB4VMWYsDULcvnWbnrwWPHebG
5SoRCNrmsxb8xQpyr9gXakD0SHWZ+YbT4FOXPgDZsNxMhmbA0Nsqi1Fpam1Pal5NOHd11VSHj6V0
v/xFXgdRBLsWpHQrL/eYejBf0n2eRvL0mI72+I+4MhKxdivuH4kyj+Iqx+BQAoOBdKP/dKirwnJF
X3hEFjsovyenRph2vyy/lJxEPIIhm6Jk8aWlAdoVci2AYcch/Qhe6BjlV2kjZGKk6ocJFL9IQPPx
YHCDR+bvfhN+69J8UGUo+A/XU42ZiQXdwy+kan3JF1sbYw6+Y9+MELLydn0LcmWnWQUAQ1KAZJXa
j3KFhWZsRo4SfuQosIfi/lZ178NzRWCovMAplQNMrvRjG+CuwREw9dPkglh03D8UgB6ftvVAO/ox
Ru7vkf+64bfjrfD7b35HraNMMNhgRIGvPt6ed/ruvKckvH/cojTIPbf+jFMSutnZ4r1jisQfcXXV
37OI5Br8MA9MFxoyUKh8INI/2bIc4Q7o3jzbEbGwKpcKpBQEj8H9TCGKpiv63Xi245W2nEogrKDe
TBQtcENNoRYLmhQ3RjZYG9P/cOlbWnnKOt0ySBnYixdGOjcoMnSFR8HGlRdTHs0RzzOtkLXkBkjP
FjxaCRAearcRp7C5zN8OzThlogwmD3poV7/CfFg9bQ8Xir3BiJMOi9fLq0ix+1zXa5J0SjmmM0AI
yT1/hprtrLUgroTN8e+dnERyJAvMieyZgByrqZOL6bsVW7u6y7LwMv0V3/dTF4uM8XLOIffXIqGE
f+NE67OVYRGdQKofGKKSm1NuvYUbeZIGXCwqqZ/ELj0w8dACqggWI1nYwXVc7CwXgA7I0V84cNr6
NZrVAQKowwcxf+7+z4xjUaVeeQEuUBC5QYfI0igdimnakWau7PoNX5WJcOwhTkgd0lxWSuiYXbY+
OyNyonWM5ilygz4dIHGJRM7ypt9fF+gLm56O0ASiaI1/b2+IP1z5BMptgnwSMvMOU9v5PIAwPSiH
0mrGbn1b89GjTtaukL2EI2iBPBSBnnluEAA8kWY6z+bZK4/Y+QShH5b7OIQ2EUYfiW9lRWktlsGA
vDFaVure3YelQgN3J97UZDaGnKLksziNBfjdd+C+pAc8cp1u8DGQzSInuAAoPWuGJENZVCXiHx/r
mc5Q9DNaWLfC5rRVc8r8bqy7/7TCZ8SHHGeHpA6TO66m+tcwUb8LR/yzrU+Vzha57BDKOl/9gh46
zyMdtWMsTF8x0wpM92e5OEBE+3eZra6bbhGsSnYrAJ3BnoJPJSK6r8pVcVMyjuem7GIUoj+8XPrC
ZjGLH8jR9cxNl7pCjKOSMYgB5PAafHe2rmMWs6b0uZc5a6VkUAnc2zYr8Ge2H6ryqsuKtazGBXSg
KgyamsATklth2XR7KkySfj2Csr3YyHXprbDlnWQYqfdBJnA5CXMLzGTqwLQGpUhMs7hd29IcYus7
nPqd7AWHkIdQrHCpYvCIG28NNY5MiYri98415wALPK9KIEjZ1nQYyuqQC9URNeWbSR0eThj/ef4w
3SVJBqc9mDPiH0r00VT5Fdj3DEE6PoLKOPWX9bV6BVVX6ob3Hz2aSo2v1Cus0S74+zngK+NfGSOk
wqNMP50KUpJCohudGrl3Fo1Nbv4e2a/NGsM0dFdZ2S6z6wMZ+St/0YRNBJwAxD6c3LH97DephJhy
OY2pR/rA2JpmroghhQya3/scRfGtE2TCEyfPL4NBRtbKWUUYpawTTOJTtL6zkHWgm2vnTb/RQs3G
yDYNAUmvWfzeEkhK7keicz8nas61vRb9zp1RBPWqhPycZH4HaTw1pseuBXAXNW2CHjssiVlReJEy
H6pa9U0k7F62nGpcdmmj8K1+k+V+Umknt6DLvZtlQq8Lzqo3WcZHG7O4zqQTGR4lWOD8DloyMpeH
lStkBR3dNCjx8X85bIL2J77WRXZY5aid6Olzh5UXasNJG7+tVWf5w4CN3oPx+YSqMXj3nPc8CxWR
hPuNjZBtr8qQBtMgad46W58yNwaAv3ycjncSr8hymYfQxYEmI228jCqXuocusrE4o/+q9BciAZNg
jcv9rKo6BrUhMrpLNastxlQP1DNTYKUMYR5Is11yaiEwvtMtaOSCMHYkF38DI3CjwR9qh2WRtLql
mPsQknweaGtZgnVpbHXC0INGdps1pgNR1JERU8t+yJ0S1gLsr0zr8EFZQ6sAX1REqXs3QRZ51qys
miQJ5QwZWrq7VnyjpYeu6292R+eWLmwja+ZW2ybfzXtwfdaE1bGCGhfDujwnkTpyhnrKCgXh3wV8
k5cOFlXJWAUdLGFhoDHcommy+njtM0gci9kexx+Ojz+9D90OVhCD3giUH+cs+gf5BQjlEKteuEUc
sDqiHcdZcKnwgYH09unrEkwWwuD4QWxpqF3UK7+AT5qA4jBXYGg0QlmxrMo9TwM9mxUTZeuzTTY4
MpdNo/ff04ZMIUt0YFcwv035ffiuxeh8JvY9z08NaBdBJ3f33V3YH7AV1x8bjLbzgX7TzVHg1rJN
lnN/0JKG+1dfpuKQ2tFeYSS9Dw/1rjJVoATzPx47O9Dhf1bsZg8S+OE9mYv4lHcrAgJUO3rJuZ1b
zLUhd3p1+r/Db8gk61NYLGtAvaSmXnGD1yedtptcrx2tGZKN6eAeMDm24JkDCqo2JsLdehYI0PzQ
SXc8qVn/Fbk2WTEoQ+i0mr7hgRS6+g4LLsHkAG9YL1MWhQdeaUv3C8uLTPwlOnYuPgRQg5rsupvv
oKwgmi5+LXpjlCp1KdmqGbUBRUt3QPQsROICeJDK/OQrUOkZ2ZMUrFyWKNUwYYssRJfFgc2SWGp5
VmH4FTRsLi3/rNXRaG+R1qsAnLafTxXaqpObW/UVtKXYKzk4IEj4BY4rj73/Fy09OuDZc1kIKle/
cUFUDZKyK7x8rORJYVXLXKJ9NlxcCa8Qmkk+MoyKQiB3fUX3RUrPQy1q0KrpYcwbPua04xG32FQG
MX3WtnyCc/Jc0d1hcygvwVvIbUoemdJjRf4J4zCdRMupFAgdOv9qb/xXOzNuepyuJ2CBEh76x9Gm
jsR+w1FQJBYpRAGrCD5PPr04s+y+9PT5Xfae71RtMOHrdJI4cZaAf9/MlmI50aJDvVdsghUqjB1n
nt6quhgY7ichDYCKMbJXAgvTgj22Vl4P/14LClYGJEyadPcZjSqC9iTS1ORgT3ce4f+VWADmMeoS
QpExLuoLeMbBjKn/Yn+BX8AWdnjUTeZQTma6Q/7oU7aj0s7CHhqriedUNPfyzsHN8g0Dm5rZhMQ8
sB8VClIlCrpuhQTf3rErnyW1lbLGs2LQQrY5tOekgDwNucAsyAAw6dDeb4XafWelqU1V2DMObJlw
tSyHNninbF0VKqYJOr0zOCllu/h+4v7hojDURRecQhTW8QatywNVFTDknkeJ/FMlXk0/OqcTTaOQ
EAzM1LnbxNPSW0SYoZ59Q8gAnO5Q+Po34vUND3yeCihthIRAgWdtTx5tke8zEdlHxehitY+gsWpb
CDiz+Q2uFLZ+Q2btZyx6vAb3EfsG9zirfTkXTPnO+lKdGQ52RIl6GrVdUN3SjKxQRqjj1GMxQJjm
AXIyMtKSeDdckuyc9RdRKxLmQiLJXnDz5jMoEPc+PE26q1fkfsGZyYlpMMcTXz8Gnx+ys93olEY0
Mv5SPM5E2MUq8gg/gh2AxC/OXFju9PvHZd2vk1Cpb+8/i8qNIKHQ4PvjnJjX5IV86aCO/LMljNSn
oohBOs4/lQm6lRYzxJars9LDTm8Eje4W8rFG3JEnAs1HnM1fyaZWCIIy1jtBNnkOXYX5nJEZFJJa
npWJiTUkDS9ZsElQF6oh6qz2RfNVMjV3WrhJRBLlApDz6QJ+gcykmzqTxwzsGdAI2ZXmZ+7gugDU
YRFGIzmrG5/tVm+QcIWyrULI/EwOTxEA1ykcEartl3zYQ0BLOOJO5iprM/c86f9lIogX8DTySOE1
hUl6cAMJ/Pg9d/bBSqkIbfwJQDE8Wb9eebuP/Sj4u+2iamk/W0JiAzV6she70Gkgn9gCwCF8K8ft
Ol74pbzVGeDAjnFfm8ad/AN9ziNFBTqLA+jLb/mq/sLxKCNK093zfb0pdNNiGUZRE5z+kLcOdYug
yUdiOJOJA2y0KRLB0wd3T2/3JW6L4Lf5saFeIAlb3tXpRUQR6+5uTycEehGBz1vTPHEViJ8aFbVQ
v18E443d7m3cDy5t3xIcB6nJpljjNO8qsWxZwlmyrqk/fIzPlc9zFP7E6x+DRNJ0hAfc8lepu9+E
qugDqhIZaqtQMG+DHSvpVgH3oGL3MO+AEMeqC3+U1ZBo7lEBADKEHlA6NNpyiTG1+pXrlFkIRUHt
SuMBZh1hlUT2BEATg+LF6fYGTckt+MN/Us8p6g6nVAbZZOMMopPFaVfBVko52FFQixvJoyzhNGxE
xJ5fmq7otPJHM4GjsuBsvDCctwAgk2ig8XSfRar5ffop3oTWrgR0tU+um6u2o5uJhw69EUhVYTcN
XvbyXtcx6AAKwOSWG0toQNgCoR8WRpZZDROrVxBB/Te7SpqvQNA1Ze9he4wQt/ai49lmCTtdh3Zt
+OhOX0UojXkFK7yJOVrHmp17I1akwlD/diS3nQp2RLYCcKpLe9keECs5CfgqkAZSgA6oahEz9N4j
p1hpxluX1KeX+yYedr/dgOvCdiPlBKZbCx8SGrSjoP5ycNDc4XtzPEvBlQIM8BaA1UqrPJSXxjFQ
waijPa+DJD9htY78NPZYWa5B9S7bCD74INUU0r62ahA7SllGdT1vBTQOIjWh+X3W2tdGrzLQpssT
2Qdo+IihrSIGJX15vqDoHL9OrKRWQM9KCqj4F/74w4ae9XKJQgEG94+9i1gWwPDiOFaZVsFHoZZQ
xiPlmq/zaqkA4f8p6Q+oWYLCkAegsvMnk/uz0Yj/ZwpNBXWMOs8IANxz64GfdmUaZnJyKx9oU8Bw
1jjQezdiLNWObSNa/9odKtIBQB/OElYtiyADRIrDIRyDorKjfv4h+g48+3P+RMby3ajBrRhqRfQv
j6r6ScVAQJP27GXx8SgnHmkHTHl5lFiSnq7qI4t6Y8hwgBvgKzu5msZOkvXa2tS13a2lRS4RdzQx
XC2+VdbKFMvxal0hmECnILlOitlpEjwy71l14sieZ6gODMHaSGQ/8AsEAezXLIzzSJU0ogD785yE
hflBc8Eja6r7tseav9Q1wOwhaAFZL6pmWzd0pSFG9aaDdNrsqGnP/vXlYg07ip4LE4LZLAxzR24j
ycxlypE2JCTw78Ty4im+tnoFZQf3ZTEZ21VkRfhtXirj+hf2MBdugsz/1bL3qqaNFuzRrKlDL1JS
JKyb7s0SBNsm4nNzBP4D9yzPPnLhn9b2WOoRuuo7SSj53UmQYCHg6q47lTCC8i5goVonzsS3CdHh
powNUScigMZXoeuBXChyXB/DubINV4ua2Z+yadsHrCvMKXoQQ1HNkQlOs0yO5C/mG5vo4ST8K5FL
nlmnNMttre2Nwj5rsX7YAIO5Ss/EqS4pdAV2vvKQaD6F0n/GJkZhvpmQHoO08gizzj/2ary88e9m
jFNf9lcsjCkkIf4O+eibUxB7+vwpOFUch5RELSQ+30pEPxtX33njQINy6fbFmZ3oTxHq/d4OI5vn
/BknW44+y6qgNiFvwOZMsSR0AfYCqsbL6BGEm2aTwSr8sTczfw4LK5jqh9+mi9B3NZQWjKaiMaFu
P9eZ/0rDQC8mYsC2C2upYG/eMKVkQ0zwoCISPCk80rKE59GFGgIIywE32j7JZi9Vqfq71BicyQ0a
JkbwYOT+uruCISja6i9g7HoX+o8Q28AhPAEn6kZvt5SoszgdtFhCqtcAtu3KXop7V8nae76LvBd1
xUU+jNeunleAppjoEWe4eWurtyNs0+9S0zb6yVEKbwCo99u4k0mo05KYR8skx2csMk9+BWsPBRrD
ndScqlvkgno2W6RKLnCjMEfvTU4BvvIozgl0rnVJKrJL4h/cDVNSzAE7a+8VAiYnWBO4ROdIFXME
czKUdZ1GhdrcY0UwBqB+cjJXgXP+L4EORCCjRRh2Yg3KqahgvuNL3Lhf/mSHw7nMy2OEG8x8lx3x
fOJt3Gaqm7+/x0v/Dskxhzheow5iGbfuVCoN2qo/2Z/ljeBUigzIA6InpFwjA3cYTvW5UC3p6bA+
4jO6HtgPhV4TCEZZmnI9npeJiNwJrb/Dco+ZG8nGXI9UW1uOscfGbtGTpAk0KNTESiCLaDV9kExL
XzuViSWaEkIaAYwyRdhyJcGFb5j32DzWVrwxOZXX8rm3kYZU+AAwA0guPKGuFf9W5ZRAg2iKphSC
oyMHfRwQMT5S2qN0cVx/4kg90bpY9qKvVuKYKdwpWxMeZsk+v9odagBly0BgtwNYaf2wLbvMhvrR
dyTxx8JPE+sZQwhru+rZO4V9/ruq9PW2m961VLy5B+8yiMnynUF3hZoo6J1VjzJ6j//oCWw4oHxT
AkvWUHkNQMcuybk614drLMvJXCkf1UurdS2o++oSO7JmWHnrX5PqXzzA5MGox51A27O9qK3Tah8Q
WGIvcNXQkxe4ov0feleifG8C1cwJinyoUhuLXy++dOmtksrPu8Paw50hrTuMqIgy322in6g/XYac
rK0/xjLNNNuzJFN7kSOdGRuoD6Y2+k056kUmpcN4ShANbWZO8V7SDXux5sZBr4DN4nPNtTuqu2LL
Aj2ivQ332SQiy9gItuEH+mChw87TydwswNW5z6Mt1jHmp6iG/b7XJGIoJFh0L2/V+w8yUugMdHkp
v4SSNMXHEf43ABJhggmG4KJCq2UGs9Ez+kg4wZ++SKvm1npAgvlhizPrzZBcdKc1pjzciZYY7cK2
z8cStFOsojfhxm8uFdlXYo5ysOckZN7gbX9fxsrnPBuNi5TOkbTMjP9q1XZLNnTpjQCRFtTz7NmO
g0VN0rod0TbURBRyZbufdR/z3mMdJNRSifyiEOpSRbIRNsM8RtbKdJ9rKEryNFXNrvxbx70CVauW
Yigd3qdaed17hARX4SQUYdSl+8IlDnILyyeKoBsSB8eMbLcGWTjeXL6xuU8Hkufg27l5TqZ7H8tS
/9K7yT+pQeKYBwlN3GSY96t8YwaEVYn5UpJ8/cr8ruS9fOtAr1GCrUy/N840yEAMdVWHEH44hlFG
B1TLEkhIWAX7tRmY/YAFnumm2JDfkucAjUbd0rYmz4z3cQtnE8fo3xzFVp/XSVCGhffHbOxbfwOX
PjzgdxoK4EMTgDYxL+aiDAEpr9rRWm4nCILsamFOfwNsCZH5VF/0FhYshXzPZU/GNVF+72/0n5DP
EKDmjmeflkOITiRvyBkfija4lTDRL4etK7PWuSOSilE+I+ynt/aG4q4pnlPsOK2kC5wDaQPqrLz2
gVFotfmRtf4buCibiVQjD+98k7k02AYFkTnFB+FWrX+yOSxwrlbk6NqyvT+/u1HbQkbbYFQuD2r/
XBsUWPFtkWiI0p8mPJSQGa8kfpMMNK9s63FpiDXkHQ+2EfSBjx1C+3iVLUkweZmp1h//ssKK7+HZ
UvRmgUustPUQWaWdV4zjzHM7rSmoUJrpFFZc8NkjlMOjVlnI/gWkxQ2r/8tFi3/jsKvoxmtvf0eT
JbEqhEWhCzbmw3uKQsAk4qT+4kUyLhecC0HxNvPGJU7wphbr/b8xh+2ImrebqO1YGMTwI5Mvym+D
6KmoO+p7TTJdG+KMIiPKqDgIdzK6iPm1HAcK3I01Gpk9kncToaeCDfDP4jWUDbO/VNDim4EqEcjU
jSifrBjRCaw0qrVW+vcWkQSgyV+HKpKdBl4r8SxvWHL/x5AKjGdEaF0RBKN+sZqYXLdnn/58XJlN
OUf93L6YZUnBYHGweTt1zp+VCssMnh20YgoIAqLZ0I0wInYiOAm6ppQhe5WwPFQCYlwu1DXo2RiF
bkPcUcMU4/is8FgvBlfj2y99XkMhwELBcr7cAu6petxV2qbhhjkgWp6kBpLmz9XbHRDIV6bseM4P
g/2+uEpk4GJsw6xbUGy4BMmbaJ/f8wlBtseWESKxFIRLoQbHLV9QnFLxS1tPqP3rupoGVQZgsDzt
I2pRDcKiExPWB5/a/qkMLBfcoM1PB/Ho8A+pF/vvwmx1dNQWCN67/FfjQhhzrHOHDMde+ybRyYIM
9kuBeUtzRDRNKSx1zvT3qx5tYcTI3RIZebEK/+M8dasu+poTslBW/LSbXBWD4wa00NvJ141BivcI
yfP6gofGXABc96PaCVV/UEpj2AyKLDYGcxRQyvE6Y7qzCXAUTwDeHPsgT+UGErqO6UVU3p8YwVvn
Polj+KMdYTihBk0lVO1EuA+P/ydmAOugoBrxfqzRoYpJFSj1U9vrjQPBD74vefDsdn19UfmO+OC4
KkEmBlpbuR2LlFQ2JQUZdVOzqTLzgTIFmc1H6Aaqvl/SaXjemslGI9V8Ib0rdxAbqhPIE/l8wiZh
4t/NcD9FAm1q5TeAZdASGgISsdpnGVr5scxajII2Rx42p/AAmSyvKNYVHdm6o4/p9UuxidahehX3
S2zv2aG3qlfATc+4P9eFkgbW1WeuPhXcouTBLVlOWzZTgnRuwRGqmyLgX2jPhlG4j4QM95cIpEwD
xrW/Cn1NLBMBzr/Q1KvwcJbcQ8XzYycV14SJyDn+Dwgdl1kV8+6dMH+IXMPv3WMnx17nrzLRjA3s
rEZSCZdIDJ7Xs3krVYXzRQKVis0GHTBrDfhcG24zmMd/brc4Sce7yv4YglQ4OK0edx9P7QQa/CAE
tO4tZ5GLwJRJswHbCydVupoYvePALnD+XhrnndDWihJUI9H9XNjYbnPEGP0wJfgL5ah0Gy9+ynlQ
WxPKb1M+SqjsL6CvnMY6ucz8UpPO+f/T/dcmw3uglGf7EX8Jx2Mn0WE9BSdKPR5BvuawTB0fsnfr
V0R+CFF+BqZqypHRFOZgzAW8fRBHkVsSKSE4ZjHrxjfg5cwHrbqvc72jGF90KOrHr3+c1UTgpDhS
4WH2gBE9ZcA+v3rVQoZs2I2ilT+oGNPwTPdE5XeJjxpzrxDxVuariIu+uC70gzI9wq3hJOt6jcUB
osv4bwRIJcggIna56fKbXJaV60bpOh0oMs83NmFjfrY9pU/VyH86XFA7fokT14os29vx6YI9siVW
WAlQmxDZ4akx2/XdO2SNJqXLFtme8iF1laiYliwXfjufX79E8wMWQXmXmWRtqzt1UTr4DIVTu1zx
oqr1aZL6Nywm22o888TMHujdtrVT1azyYq63RwLmN+bdZAENywdxhdGXYsIwkQpfceQnznf+LpiN
3u4WXXGTglA4eoooqSC/8umHftf1x82ej6DrbR3q/bTHfYEJvrOKFfRGiFd07LM+LCgUR7nfQl/n
WnSCfJOlIHBp1eHhmDNz7b2XEMO7mis/oMN4HzSBqi1stnauKTYhqmnK5YH3qTCEttzhydJu8hP3
8v9XjCWN1lNEJG4EO+cJJkJ1ags08DJZOzbX4LTCret98Wg0+ghkkavVBgctS4UAYbUho5Y49GTG
i/6ONjI7xosPvU7my57a8IAv+k+pyUXWCyzQ8AsH03RjsHw+vpBgKxd8mWajaT6uQKtFUYe3ghmv
/3zJLJlTLOn2MQgrd+LvsQad43/jlFdacNXsGXQR61u1BWbDK1xawYrdIeJzfWjczyyayA8joImP
w1Zhm6as80zzUeaTBYEISsW8fwtB/7OPTpOk8RnsWkL/u1pfAcOXCDo4VoT1OytQJsAtKhto6ahl
zrIodt18IRDcWsVJEu1BEd+BCA2aGsOnyZkFAZNiRKB7FFNRSKpoY9DnTaSLJZLziE8bjRNKkE9u
qQwWGuqXQaf3tP7wCzbSEvYY0AkwfM6xQ7LcQNJ9SKh9EYZ4zV9r+5nMpWtJLmdwdLtekqOEVnmN
TaE521gNi/CPy/LMGmvcTli177d64X0CTpeAth+XZwDvKEwqZbXoCYPezjWs+zGN1mvqUNSqx6YQ
tNnnezZu4uxCnFPqTpI3upSNrYOgJM8XxbhF2tf/uB0uvkFY7D4ehsfLY51K8FFCDglKk9jnOPu2
sHpUIuZgIM46ywsd0emhHgIfO4Px0Tz/iRTql5eNbcY7CubNCZcUzyG/bscaIgl3y32rW/8EJbdl
+AF9KdxFnlJsmNfVtfQl5WrGxw6DRrsSYfae4Rx7LUcImWSSVSzKMxCPtWWBdGzZJDN69Q7yfwN1
/NaUyGBYNn0d98CAck1y+wDww+gxhu6UdNnnvfs9KUWHpvqPOUah9n9L4VxLOANF4ykSinT+qGhF
uBZ0EGcIs2Zkn4qqHo7BoJsO3bRYtQuTIkkj1RRqAfvCEa2u6pdG2rEpEYZA/18FTtjSzVWPm44B
61GRksvjqmF8MD6oCuVRzgomwkxA1rFfHd+Cdnb8qO9E8Pq8ZF6h2pUd8weKBF33r0Z+ljdHFkLg
YVmI9w59zA4Av78DUB3Vf13QpiK431NfLO7zzAQyINrParHQ+OHv9lB278L3pYIb5XPozSgIS8KT
X7A78lYE2hGn09GXEoAer3VrOkxB3xg0BTDemZnr0kKVUxlejPRZpTkmFOtUsAMImPvog8fuHE9n
O22z1ojYkxc3Z2ksM+kZb0fzaVxGoIcG7TXKUTZnBj3HhGfvKowo3Fr8ODuWuGLXgHVIK0rJ5Ztr
lcCK/Qno8iMF8KPRdUg/tuj3LeqRhZofrb3ug7cF79ArveoDfxzIwIxqkshbInqEL96BvMbbpGKo
q8K4h0pg8Ykj+D5/A7OZrpqp79OS0PfrLdtpB5U2wTjNm3tFssjVvuaICdwaNGfDcEh8Ipq1ZD++
qvtyLtbyeLVLFJ9rBW2HmFfprJicXZ1d/R/r8nyJW3+3KzDDjE4M4ADOStlWIbB2fARrZOqXGnCK
idKbPeGNkcp+WDSCjpXNUu1QwYgnywYR1XpnGkpCsh2M0bgRDNdZLQ3Rqws3SbmXo53zZx7G23bk
Rqk04YgPitlHP31ddnWfqmnPr/LAfppBFHYNnVwkpy+24Ejx8eMLnKnRP+q8ijNS7GT2aoEZ+jbl
eyUy1O2xoIYfkaVfvrT4PnEW9F5vE6ci1fl/U36eD2GmJB8tmL1WDF3zEFbRBitt6onfNz0jfnc8
j7B1Omfe7UDXj/P8CZP+N2x+3LIro4ODl9Wr+FQNVwnHNVvK2QdkOa6TmY4xaQsYCr/h/aW5PjbF
LfmX+mv371gMANF8Q4K05UuDmNW9IxgCzhrafkz0Qug3wsKmP+n9WhfWFVdpGz6kI6fcaUYXZMmw
XhN/vyzsNcZlv1zLHT08ULir4wBUl9UctSVUExnjznbunox3KmTk2ja89s365PseRnMAvJkc5WKC
QFJmXldR+AkVCSLY90ciBquxJ8h5Ak7HmLlZAuJIFRVEeIsplIKtHkY2bG7MbiVKQkFBoKg+oON/
75T8TkksSudQl7hg6X+rS5OChs33Cggw6icDaM3YlU8JFVOa9GGweXPBCp9wSe6Mbfzhrctsy6ce
W2/YeDTaTyc3qgCERfUEQXP2v19SumD1h/gJtpsm7Czjyq4Td5k57/IMbfMSsEw1mhZR/4yU1vQs
W9Ei3gkH252QH+ObFUk9pP4EhV9t1ZlEkZtCbV8FBQlhP06ka6y6zDWWdt/ojor2Mb0WjBXdXF5a
xOC9AqHuDbUDtCwh3jcp8T2nlPtJrett02pocButkfMszQt77R5Kfz95rAf/lIT0TRLxBbmp87MS
ZaOgENEDgPWf7TRuYQ9XqNlNMQQnh/KaQ9ETQM+tBrvodCcAm1Qm4OolHqajoxOrLgh3kUPaNyFz
zMGU+Q6oii7G1IweDamx7nUUMx+WSJgyBEPfnkPk4j8e/5F2qbrO+gTDgFwX8BJyaYpu65U8i3cZ
3Tb9OJbbKAODWpZVRg0h0Aezo3KAc0L7iprtlUETSJyyQUWK3YYfPQ1P9GlJpXRTsmEeS0CpEqHq
SXwNYQgzTOmaq0jD9p+yyaKOoYTApNU3rsDIfa76HLPacjPBnDahpssyVZ6Qrh8TuhFts15bRVPq
grZ70RsGp9Jt+s7E2z+Kbqx37xuzeaePgwQoKWtRnpHmJobBjCiOg97Cgo4HXj1g/IOBw50tyKeI
vQwxScQNIUY39WKnFmS43VpMDcSIdxNxOqaZJ5/+OmCGm7uiCLrEtmm2aN1nqoFVRLfiGD5TWz5c
cCreLsxGqqtxcokGkOnCLMjESmYFViSMCEb+WePC1yRLkwyDK0e30GJfaPM4K9hckL+LsBo3WhCG
0Bc0J5ISVcnR9HAu822etj8NRN9B/fO6rcHkKjTLqLAjQeWgBQf/WLKKBgnxVDGC+Ch5hVi6LL+J
d4vzm5np3s7IWqXUXKONTlukGy3q1JjkM2QCiszJjZ/k4XlvVRGheJEftSvLb881K6axDIKmdEyG
Gv3ueSmBIc+0DtzMkfH0e7LRz7qhRIkyPW95WtzO4irUVhbdHFUfGkrepj0snspn11IfRuSXw5vQ
tv6dzsBBS8o+ATLzjgItkK5vShTyJuZHRJnINVQxwbanhfgCnmoscsbhup/nLOF89Ft4Py1jSPF9
ym48SdLjgv7G2MbJhE4fIKgKekFnUEv0+9oFMpffXWs5Gp4/MqXBoex4M9xWxt2pgNJdp+/M+qxA
jFFqczzCN8MAHMqxOT+4mj5y9d25SvGvQTJzZe3T6aFikur7+tatTzoDOpVUQtvKeZKW16RM7JWn
QvvUX8HEf4ldwE+Exm8I0IHj0ikFfKFyZRZJbqH+WJQUGy4smvX0Rssa+iuun52MxOKE/wPOXu17
1ZkANlzbFtwAP7BP2q67hdKcSBIH8qdFgEAZIFhTAb6hBNGup+U+3qILcJPBNLsfTI0jSHB/HT4v
2+IkIiHei63lwD01hzBmxv3LcoIg3sv7qpd5/jz2SEeJ0CUo7MurlrOX2xrYcSfTQtM+1Zwv5JP1
dFimlXpzlFvew33M0yBY0/na2mCaOKN8xQYGV0nTJQb4RhSdCH3+p3T5EqyF+i+71vVNP/mPPtAi
ZRB2bKxd/DurQXZ8YfpQBgQ7JNSnbKR/ddfnOGOwPb3LgpiIyhAKxre42H3blwO+K6RNks+lGil0
6zSHMlKeqKYwXiYF0nSozFuOd6vFjrAzuNxt9ZvUtbSADr7L8QTvL4fm2Zs9B+0ReE5m07ao9CkF
bGiaDMBKRfyf2lEFPzh76ZoTXh63OKdeOHMye4HQSCp0wJbzCywvfkFrMRyzxvLAppAKWdfNmfVN
8FPe4+S+nF7OzRTbkiLWnE88TJtODsCT9LcaZcYyCdC91Tc+H0emMH8yIIAjWGy/YS54Td6pgEjP
HNe5Fu6wYqZYh/xSwd5VSp4FupvWOg1gD9NUkyPWGBYMiVIsqaFzEo271+fUf7aT4vSk9h1xRJyS
pbVdJv8F+QTWFtCYf+dpfOa2EM+jfn/HHkI1sDp0Y2R8qdOXf5e8ceAvCD3YHeCUpH/TQekRGGNm
2ESSVewY0cESGnX3+hYFawh3y9aDLyQDaBOv6nVkow64KRNymttpX0WYuF5IgolVLVzhd/0cTkbC
9HsSK+9wW+PV4zO4f6aYE4eaw77OZWbM/pv6xPyX8f6H3LuC28oFnDxE5Ga5amPTyw6lTnm8TFW/
01fJNujgcBX/IgLwtT52heSFp1wE7f0+/Ozlqt9gfjDJPD4oYdCbrA5R5cyndsKK7z03VITy57tt
HC46ENXw1lObx7QyAnfhuIcI5Gk8wpJWOhQwDP/4+/BYZanwATZq2+FQUH8scH/kkpQ5AUNepP24
R5PULYOlqnaoNAFGdU/qpcf5C8XW2+DVqHNufW5C8bLdO91vPrPiYCtEoTU3+Su5XcEbpNh1luOp
Fe2IRH/5+WOsw5vmaewDKkSb3++0MZSA9VCJShvhSrAKl68Nkd1s38jX+R+l+i2w/6YEiVNjTU29
1spbAOrt8CWTCjVzAHxpRCKwwk4jsBcGy5ioLwNHqQb0K0pZIPmyRu7bbXQvq/8/y73iKnsBNztj
f2LpZsHrdyHnwPkw8UWMpTNFixShRI5wN+lgtg4fKP6fGdchgDb+lsrV+XYWGbA6pL2mxE2wED8x
g1tFrC9ci4G6irY4uul091JJVRDZ5ZOVpSwJ1JDyel8gz58S+uF5xFMEPAYTlVzhrdiBAhQCqEeH
yPHlrkH/Affz3hs+3TV5ew/yIlUVaxFmD5le9ufCfAwjq+TnphVshjDp6cIQEjf+SVd9bWVK1l35
ULOPS3Eln9ihEA0UEW6ObCmcV8+lk2cSbXU94AhsBoe9duWJGJrR1YjUjg3majQrVA/HK1jjpIS+
B/hd2NCDcJgq2AhqJmO+NN4vtG2KV6khy6dsvUlQwZ3mEziEZ6lkV7RSke+RPkI05Nn0IF8/auJr
JGQPIAX9rLWkY30FfMzAMgaExC4aGZC2LYkbuQ4NOdT2BgXQWgaum2MeXNju9Ng65QopxoTRc3nM
5o2XAGt9C444Xxv4IRYONFT/hv0KS47G8Uv8n0IQZGVTMeMTRdI7z0teEBTLhyyN1Gga25k+NcCm
tBb6IqN02s7dc2nZY0XmKJ2B6Z2tn7/9f2/GNYrCz/7IcnHu6niWMTdzQjKHXSHGo+ZjKR9qu60g
pCCWWEya5ww8zVoz8HhV846QHI9TmCoDCt06bvfHiyP+EtzlTe4+xge8XmhpwZmOOBYbeVuvlCgD
xkeaTbld5QFM7pip6WWODYKytXgSNf84s5zWVJdaRmpRxZlDdm83MPQMttpKs1PPs5kMtX+8NZjL
A/ZniJSCz1sNoAqCMLzX2L/JsaiO0oeU672U0mQhs0ZQ1vXYlYPZqbz3At1O5WO39ZVHkWkKKjBw
VAsKMQDNrl/GA/2f9bqTG5vunTbUCyd1IyDI7++HazIoH3PJMdVmKzzwdyA0xcoEEfJG6Y25y3Jv
FNNwXbtRTJMaTRspEoOnjrMN2Z9Hl+0zSuNDJ5BxykF6asRB1SgWiHg4Mj1//+d3bGk2KgFtYfpM
SZ1FE7Ssy/4mQ6cHkaHdJNldZFgAZJpOm4OD9hEXyH5gWRcbWnSRgw7fWhoUpK8TEGfOC1E82rmc
Xjqlh9dapj4H1r2utZoiZr9RTLd0YeUBsmY5jD5Swp+JZhVzagunKJ13g5HnMVAHDU4LbP6C/rjc
j4orJszWUf26dO1Sdupw5K7Zw1e8rBcwuCjx1OgNOJl6EaF/67ojTcH/U7Uo5kgV3Gj5QHLgEt8W
JEdkB8KJzNEDPOIWrutj9h93jkfT9WgLPPRvkGPRZ45fVGFp6GceriXiX75uIRDoa+Y9aUjH/1m5
hK31BrHiqY4HohzZZuzvUx8HpxU48/8AFfgqv6T8Ch1z2gOmI1cwAhqmlv9xtop2AULim6beP1y1
J5cimCc17t09GY93g/20TceRuO+YdErK/VTK0Bnt/V5PnRXFIqXyibsgCEudKfwSJX53e9MX0FGf
XywpZ48lH00YGDL8VwnxlLMhUUNvCU/PREVKQHBCF/Wv5s+YhYPr5M23HdI3DIGPJPsmiYcRnizG
UpiGDrfuFspFz8NEorEwDfFC6l9O31Y3OnxvL08pHaCw3hwvcm2BBI8soNXAAva+gUVcrm+RwM1Y
4pXe3XNIllIC4hVfpbvkAUqWQaLIFAndXQFWwSIEA1wwMqUTybajiJ7zOHeyTp2MCrx3rtiy9HDz
SlWFkSMV6UZ2FHnywZfAe3CFfrYtAHdLysiyQ8OSJu7HrIzmpEObBzHYVdKo8w8XSlQnlE8ZuxKX
uI56p6pmND18bsk//9PLYXEPuZpMDumtZfx0HbJSERZozFtjcHh1fbGI2H4miY6JKVZtIvNF9fjy
eGzkSIQx7vXMxBJV6ednHZ8EgwDLkjEh1DUUBmFPg75M+28aGfG24ysbejGTMwPfR0xZ3Qr/ilnU
5Im1CMv+0S4XG6ujsp3cc7KfqB1vGKwnLXvzKR45HVY11cCZ4hH7WaBnsJRKoHDI8RyQaL1sff2J
joDVH/ETNGxM9QgkvUJ8hivVem5juhuitGnZJR4utjNpx41U1dEwS4XmNG+g1CeDtSzdP54iE1C9
MVV5x75iU8+UUUG0OYY1f5QJBsrTGXLS7vrcy9nTgsXLPQykMrwe5F/aLE/f+YMTG0A33+f3BTHU
/sjSSbW/4umLlL8qcP9ERNH4mAXTBYyR/UUMOw58PGHqyKwIwJAWzNmkmkA8lrspvb5YRXSL2hUV
Z7RzmM78C0/HR7/rVWRvoJPZZOjjJqSOpmD6Hw3BNE/s+nzVeLilBYJviyxUa9KmucVxV6YNIWsV
E4BvVGgnLIXsscoi7m6iDHkbNsR8BkobM5ECzKyjsOg3Nir67kbgryMa5YpKTs3rE/diMbeSEBth
LHhWZS14clXp7ywRQ7Ox7W4vrMSnpDD3AjWbXBcLR8pfc99a0qLFplizoS9kDN9ewa/7pG/QHetc
g+xizWbQcKa9Se07cFeILL+B3jxp1vxWfveurKyIEJwgfisH2CJr2yd27vF85GxamsDFXZhjqz9U
OA3HT/XhOQFU9wcC8d60U3TQv6Sd8qKGv/1tRJKrkS/Wb4IUvuhX20aKx08nSGqu69R2rxZ+0T66
XL46jwJqYTkUJI2fQ4B2fcLaHx+ChDmT/7GrppsjrdepNBbQpdCGWIrocJmyxWWW2/lpMINE8Xlp
kMXzGgFxxyQYTkAcscbx+AboLitG+iIdr2PvFFK4nrpNc3+r+9pTi0q6gIitXrtPkTpY4+zKA3OQ
dIRpWY1W03FZ9tQ76qpIgADENi5qVbEDyJvPLhuNCkfxwhdaemdPcNZXlfRWQIzuwA6UDTjJhCOz
YKIWFXb4Aft4zXdW0GPtKLpqzaIS1rlV3AMciHepsAPzKEmP8exlju0OIeeGgxnL4vRS76DU525o
4OkFLCETC8ZECcf1QqzfgARReWzaQkQfcvJ1XuSdE6MGUmjrtUUnorM/FnJPI9RsAFyV4PcPopbe
/dwjMlTkRej6nsS3t8SoQSJ+7jtW9/WJySWwlSxzchMVtQBzV+YYRkOKEeultCnPXdg/yCDgg7t9
jW7xZyv6RfXKnv9PNeSWLmYxl37fesYZu+nNm5zzc+MhFVsvPNfa+dJxIMAoCM+UDYVTRT8mW/XL
DM56+jgqe9vSH0bgP+gqtUTXOKQYjJgg9ASx5KervXNf7r83ccebKdN7RUnhlrUwdAeh7Hhce/1m
pSBOgQ3FgCf1iZzf71Fdts527WqWBqZOhpYuZRiEo95/xpB1x13sOx5yMAZF/m6VXnF1/IAMv2u/
tna3erNf+h1+5LM1K98yLsxmNOBUumWSoKdRzuCEq7asx6IBIgzuBdgO4adnMia/aI/kMrdPa+LQ
ki2pR7ld9NLrk1qtpw4HOTtfmjxLvdOJpqNuepoeISSaPpOqLEfzwFZBV+ATd+sK4ASA+xcyDoZZ
V/ynsjOoCh3Whx9HgRkvHgC9ZXty34c1cE57xaOEQ1uxSxe3cSPnYcu+XRcCgYO3d2iZuL2TZGGG
JcWkNjXEJjldoMNlK9Y3liyX32HNmLTOIc7Gnn8fjH1rzZPwU8zGplLT9Aa5p+d87dZQhv8Oaoi8
n0qcdBVKhV2gQU9UICBkysqCB2LD0SWIKwq5zw0T7AF3ARupmy4YZxTWu5yyxIysSyW1MKAQMqiL
y4rZEguOVjHpZGMheqkIthyuBud7a2oY9aj3uL4JT9H8BfwuR/x35SBn8tdFvmtL/PXZdeDjbSKv
q5XPhIdEGVv+ViXirCzZJyo+GHdFaN7IB29o7GetANS84bWlSJNbNA05t2f2e5FR2eWdage5GNwO
Nv0zwtnR5/6Qhg331Urvu4ofDpfTV38yXis5KjGQxZ5H+/fYP/cH4EmM1rXHN34fi4fPx0/hUkq8
l+VpWuRMWXOJfcTqo+5nd6QD8uBw6bKNHtsEFDJ06raMZDd4rq5KmRuxPzDDh85llzJ7aW2JeKpJ
cAeHuuhtzr8gEc+E0/QDvMBU1a2cvbsrox26ceLbY1Id2zPHiNVlrOZcPhgEL44d+exZJohptH9L
Tq4fcyhZBzaagrLwzkDrV9dhKrdNkx7gSKXtVztHd0XvBwjrCg4u+0Pxbaf8PXlkJg8JFxzgF8/p
tmXPWsZCREwFHZEvy6lGkYOS0QsY/onfZEtXt4Fk+CxiHjH1WRfO0b5AZq38uk9P4Dg3ATS3ony8
zmGWVOZDPg0Xy5w1Upnxm90B1vy2IFN9YCB+uVQ6Ck38cuUDKa+4wyJNV8brfHGX1fhFXO+wt6+T
Vrz3DU+ofZp2D0KKTEry70yTfVEyJllVsH4gsb8nI76MMZoFdiij28hnymsRDqxDR9MsuNJD/o4Q
MrJa1qk7vDttXDB3SwsVvi5t1Xt6lKjt9mrK39qnfjS0bzhTDxtWCWgAoU0BLLT1L0IzoXFzpDbf
2Q2Xqz/CP98e1ogmd8YA2BZiStv6sIMVgbtrsBGcP/2qTekUI9Irl/aucchiOaMEwEwJ+9pvUqy1
Kj7csLMfgwRhIhR5SMyaQqhK0ImwrW6JnpsBQuuxfxeswmhVFZFhu3KoHAp/uyNnJUZyhwg9xftS
PMNoihciyCBKrTeiEv+DPkNiRuApoMDqVj8ytf2zvpY+M5Wv4dqNVUSPeboWkObDqoK7DNS/0VUp
pHpBIOLTvIFa9LwV7qAwE19i0DF39xZy12UIzMw+HKnW7S2jy7tVAcdxhHw1LSrMKn2DxD+08JGd
uKxdl7KskFySoD6JEyWeGIlSGXfgXv3Lx1VwzqhYJNGKCnfy4WGucUGdRfHeJH45AiqBHSj3p816
ER3bF4akmXr7OXd8fmYfr1+lFwKG84iaieaJk6sKYfkrMnN5l0xR50BvbJiSn0gTAAa5BRSHtv9w
uSnZ3pXRpG8dw146l35cThtcH5Uut6bXFD1d8Svwgwtz5H1a1Tl4dZLKbu5Sx6Qoc5qgYYtQ431d
nqbNYME8PxrG19iqXl8B66mt2BtjlEt8MORva1ypxrkt6szXAgbS7BzmJkEzteTuVNowLQla7F2o
bAoD3sDglRs5tT3bpMcsc8hemSSTUwDsnCokfHBjHUDCS0ZSjjARclaso5gnXTB1LYslib+8FyOt
0NIbO11SrFnfPT7S6TT3M8NLTkwuDM17l2hve170ymalNYcdYMhZBcXd24KsYf3pJUaEtXOksAbm
oIUOV5KTkhP4qx70Qe3l6wGIMZcD9srE4qjYOTXmq9kPOJwIujuuYP/nIVVf1nEccFakHssw+nYJ
IsZXq3YyamFVuhuig0ztselTxbWNIRdDgbHlm4BSn4B90NX0/Lr43kW6iPUpL9OEnIdR4nKzI/BZ
FJ2rHjjbilG9RcEU/j3ZbrjFBqMHZ7NBxZ2bGjKmjQLltp0m4DzzxD3Mtp+e6nAZCEPme1/0NPRx
lvdEtP/h22lk0+/CI8HBDXHjpRKtTnDlJxpQU3IvV7ywDQupaHrtxBAbQ1fyBk/YOXg2EUTSYfaU
3V2V1Ddf5q4VyvpuYFBMQ4F8GxyyrWD5/rsMP+YsdlFdYcKYN4dS6v5qO0D+rP5+5+l9/DCVQfUF
NBXHIqDngh6GhdJg9ZN3kdA1lApT7u78nu3+iMXEMt+5hgBuepDO0joAewC9Yl8fXrxRW1aTHQ9W
uATqtlhsaJgXvvlqDuPkrHztWD4n1afShchRRDdX7UZc1rRCtjRuJw+G90coH2sxVhx43YqIucak
D16k6PWwGQJWP4W8zgWi45YpyH1Z03HbFE/Vru/gouGrqsFpk6DBF54ooHnukxagNziBrHjwI69A
dRrLaiT7JkhY7uOHtKJtLD65FIb3PzGAS2YbLfDe7DQhLGKfFooLz1J6xo5JPdc9dBWhHWLDogDu
SkqYWE+POT7+3NUCUBSAHMTsOYJ2JBhn7mIn6qsuv4TNTY98iUbcAsH/Hj3sc4dldSbuULNa10tM
BVTkL/YQHIgju3/WQKaFXlljDIb/HSVK0tkZ/uh1UDeyhHfwGnqB2V+gCpKWw6OC0bm9bviokyau
Cbl8m1V89OKsL+IncykmjD2BcC0f0fUgKH1gWF/HP/QW4rx/GyFgOYGF2ycPgcELZ29AnFj9xH66
ccckGkdTxLLSCuVeFMUhNWjvizsQXHIuqRRIRNM8fzAG9yMnh6gehPGgDDtUWl0KGDHotifi1pjR
sckDleYAb0C5epwrSwIfSA+vvdHGvGDLQnkSG2P+BQupacrhd0ticIBYNRWq1oAb6FE53CbmmSMh
QCTSTWTIO1G4hzZBYuc3Lwc9+jfuOZYM80lsWZ3YYC7nH+WeqcFyuEb5C6+MwznUkkrBlIISC8C0
MFkZt1YwikeGDurmWfGTKfedtD4BlGNHJ1E47/VswMn2XrJDYHajFdce2Kr0RZMgah7reTxjQqzo
JZaG5iSZGe5iM3gtiveCSfOdokBbQAn/yFeNxmAmqBnxPObZtpvqg56DTsYEmcqabLk+wztR4ehb
s5WI0oRklz/HTEO6TZVfQpoG0eQxlhpYkGBAC/oEsP9GKQ06GWQ4qzJqzCiqaz+/jqxAjCnxMjYT
4t5EIGd8hpe5KjIAtM8ktHAkuymTKRx1VIjyM5XAosiVQeTVtx3xOkg+bJNXpK7lYF+ZIdoWywiD
coZkW3W6GfR0T3I4Gdwu7c0XUifQd3W6zC7+kTr4u35sbWkRwu66/6OoWn3gdR9l7jNI90EngxeM
qkj8PSKm6ljUg2PHmB5mIlPocKikzDD27cg2GEBE9Fd2vpDRVnrZZjdhx2sedRfcllu4bcUzFpdF
r9FjMbVzvRPBToZ1ee2VbrjkSzZ9qGmfv1a/VArmyjn+IUMLYL7tUu0ZQliv/1PN2wktSjT8/rjP
ujwGIAWkzI3vO4YJ6FNRVlCYHHwAX2jGJOxvpQdJliDjKT3UpQhsfKqD6YkCIAneCmAKXMQ/c15x
JXxINjzs3zS01ii51dVuemLSIb6bR0SuyIPwJ9ero8hl/tQcaRzDOvbj01y7CxfM99rJywW8fp4L
pod2u1jVSD6w9AaXWGJPz8TY8gvKImUxw9ota1wEFW74Ci6a3h1nVzFR/y0svSGg2ZYt93XMMz5l
3YFsC+M0OLVUpwRcKvJyqDF+Mvh1ywQPyfFpYNsGcbNLxcgQ52Pn2dL2w+CZ9x7CVX63wIGVVdxb
AzoEb7SlDF+mZ257lf33+nTZXozU22CXty/FN4G4SrEQnvBeebBo6Qy0TqtDl+4qVpSPCL3T0AvA
DyUmv4TRjd3FSioeQN0WUwan96MBADopCwLLeN8FfAgXT6sZ6s5KVdeYvo/92glIKrSspxdmwQ2L
/2hZ3FndVEiA59jHHZN3n1cbMyBF3CUcbCC6GFiCX1fFKmsC6X5yhHF3UWj9jC33jzDVKYj+lmxg
j9RffvanBqqahGl1MXi2SPAGuqcybmzpVF/bJvLBD5S0ezUnyWYexNVqTycrPHEDs3wCTybLHGrW
K+bRl2ub28saz0hZ6wni4/fBkL262o24v6Xgs0oCZLEWLcIWG0KVQ07gwcwhEDc/S1Ul1Ap6zUHi
FQoZomfqPiwMRGqNt6lJi2Vt5TH746cwA38NBHfU4ULtuwFG2flobVndkGOG6O/K+hSXdU4wReph
hZyy3jSPRSYMX9uxrRFDZHHWhjy9pQHdvqD4/b5i9umE1iCcxPWboaR/dsBKM3gT9YH1WyAy//7t
aAnHKueG3SfJsVC4NPy0hC5JpHpJD0JoEKY7zmZmwIdlt42CF82wTLQhpOku5dkZs0eNqw1S2LXy
aSrMt4EHGn+CEIIvoezRmsQTkMse2iKg5s1yhHGi9KHPvu7iP1WqakCeG7MKA8BiL1vUNWIIrh0J
a01yhHsCflH2Px9jDlC1P/pmhsWclQmIRXXLNDD72AQRVTwYBM7gYPibIFSSFLC/YrqoN/qcvflk
LgUqaCXy7XuYgHLrlTdILkUV2R+1uOG+j/jx2r9yohkEkyrpuw326E4Tg5pqlumYaIYjhMjmW3Us
mdvmLUFY2XtmIkj3F7kpNAUcYyD5E5zu0o9Y8gH4HO5SVy7+0uEhwh5+dRQp0/p+XpJ6m+2doqhG
BrxJ0cgcmZZvQKGfZ4gcQlMguwNdaBkKCYb5/RpRp7VzZIA8av+U2z4ZSMzH+A7tMo0JOprNl423
Nnvl0cJfUFDj8e43DIltMaUo9wQQyONcKWhd8X1wHuNTZmxKTVHw4eC89P/15+YuIxHmPmMQ9hh9
rRzr49HybxSH9q6allWAjFi0hsGb7BQ2xdSf2n6WaegFmUerL6YB/zwLpRRg3so/75hd2pkQhiDI
GR+tyu8JcQun45ypa9ITe52gKL+xz7ULJlqS2+yfNUXQ1nyKn/6udGmRenue1yYmsAWbrd4g+hNo
w/FOI9t2dGVgKgFmCmDBQ5pltA95Asob4npWwLVidznm2HQpN2fn4NpmHnDt0LQG2/b+XFmc/qQe
RMTk5gCFyUXs1JkTHs9fO96bEsY/6T/rWkx3rBrrpllFcp41sWOj1d9gjkbvvFhM24LXVA0qnncq
onV0Bi2ka+MXJSqEFp6wIhploBr4YygaVO2JExxz011FyO7VZNiO5wWgG84rSnlRgOM34t/VW/n8
1jX+kr93JqK3/gHzvHEgvWxFblLgFR9OsJLMmljDYVSpdAL/4kU+FhfugQqDNcrQwTlxUaFh4Xmb
mX9lcde+iQNpUy0a7tBG5jzF/hFUpB39kCl8sHE785OVeVf4xvsWXnFyHBICR50U1tiGbGNlfJme
rExswnatKKXM0GigkxpulQqiB5r3e+XycmafW/2yA75p5HwuC5WbHFXhxfmudAm3unghoNW6suhx
VobkyR+gjj5CHSMxL+Q7gi9T0+odFM7AI/l/AczqA8saO4Mxm3JM0oygwnde9+mPHOnBtiLHW45k
SgMaj6BxIvdPGD66GwBwzj9CLGsOKTiUMKf6ArlR6a6bIqwZaxTkCN9HBtnJD69oFMYVDzy1zotj
AK/658LW4oQtmrgLGCh88+KFnWqan9nfMSbz5NROraUrq9SenJ0wXj5+xcTgNJ5YsvY26jasfAaj
7JwGEQETEWOcYY6j0N7vAI0/oRqKSgsD2OmPs35fMru35FVnDzl1xXv8qPrdyOGWYJqrGWx5X9Gv
7ZtDzOBM8TxQUmEUTMnI6uSCKCLz9xHEnDY3UKGUbG4otxtY4TbbBNWsF4LgG6N1FPndD20kQAjf
++L2d+pkx2+AvMWM/ZPaKDguEP37HBYj/t4Bz8u/a8LY0FuF71WoacRIlYrKkAD97nlj47ka7pFp
6DlyvD0u5bOupjm4PKa3QOTa9Ki8YQQLMl39JLJxOHuy0dfZczqKt3/g1Ik96t2eY49fIfvqaReV
kHKyg38ZZKzMs6E7kWPa/DEv1sM15yYL5vnKesxg3qYyYn8jgEXaZnBl5dDLI2IchTnqOs4IFECS
t9M22Du2MIDk7s/WLC2bQI+FQM9JKGjZs999qyxiRnznGCyt9bpldGEm3YU5Pm3pfQe+7/l6Cy2v
iD+zoo95QEvRM2FZAOEg5yY8znQZa5nsgfkHt6jJf7PYzHBHvn669vSM1gR8fZQdIVu/3a4X3ct4
FUM6l3+kB5JtVVA6/IN13zpCnQ8MIbx20hPo4vwKogDWheQIlNBYD30xJ4zbF3hEFhaOykVJ2xBq
XslMhfhv0kkml49AhWKgaOzqv3V//yzckTbUsYJWu7wPZe66UjJKQD1He2f/G49txYcs3Cburcbr
1q45bk8UMHJ1cDHPjADfXLZHz9Gpa8O5yd2l9jvgfgZMdDcbFYeoJYgzqLHQApVYCeduHmPNQvT5
9VpcdD+Mmi0lOp/a1kCe89Uvira+jQejTXUvmSO0oD9Jlrn11KXH9rFGkC67BpcSLglCHn12zIVX
e2/CqiwV8c1GExR8THGlfERnhWN0dW2PuyXYUoqjjtR8Nt0+Nf5DYVjYvnZs4ObYM+jgxYlP2787
tJUT5V9bURdQ8x2ucA3xgVqJudOxUgOLBBL2kDp1uV8xPXUvdGX76Ly3+o3Lmn3lOT4POGG3ZsAN
2czO6tCz0CgGzrnqNxNJEFMwb/Zib1MZ7Kx0oOngRZp7LV7VOKHZNvj8Ji55MBoAPxjJPXm37pnR
XeCyE6TlkmaDMTKvwNUMBN0a20FuWgAolfRiwT4gw8XTYpihHfWK+uhalxJLl0TCO8RueFIzZjko
E0Hr201pQ4T89IQAyVkbZKsrtZUnt+Pl/g5z6QWinMBcJd9Agr7QpAWcDzVdSgO0i1sFWhFwHSIt
mcGRp7tGHrxgZwY6ILRen7LEj690sTslb9Knti63KY3kw/RGEAAvomDS2/ApG/UTEPnI8trVcF8/
fXAP6uej4leTpOYCGVyvRpe8l967pKaOWgdfawOTVoP89A1fazOLUjOjDXvi1wA4JbAmAZBTnm1m
gXsJBYeoqB9LbXyM6AJ+8UUJJIB/BZNihk1E6tzDVimNUJEmCvCJQXufoDEUSY6iSjdAXgXXkN6s
CzIWVLQmquW9j3ySFG1YPIQNyphXdfMyMTXCEaxQwKE86UyRc8n/tHDVMjdfzisoz6YNlkEjPyFy
NuhhS+SC4T0hiTTej95wz6eitbLO0y2rubOduY0qcAoKpjCyvsjJBjZGu3XfbtQsEa5ZODUZGdUA
zWMw6HonTPpeHbUkycFD8qx4kRstotB7nuz4y7iIrRbzyxFpCSlkgVEwprbKBu6kz4fIKV9IkE4Q
qNOUUJY9ltLkxT+trunBXvm418Mv9FI/dJEzioC5XPAD1z+vbFrD0cpD5SjdQbVWMIMWbr24MVIw
1QBY/Gi/L7WjaSLJLw8bKS6cQS1/8qJRf0Y0CjR40FanZtbu+GzTx5btMyQ9SJ3ipg10cUwcbrBB
yCfdQB0braBSdLmxGhu8FTUxBOJ/w90lq8kenZz0K0VosqP99+58GyjKlyZj9Vx2/1OAN3qP/WWL
5+o30VpZflWxUb8mxMVyn6IRArMz3VG/8BLSMckMpCZHVWs5So3FZS4M83er+ZCKqnEiTpMhFd+I
wwDnC7zqx22qyRgtPq+n+nrC6sxD58ycPzIeAPudibnahUNSL7EpfZELzwhYRsRGtkdHYb+bEgy/
G1BnHcr2gXfwBQlmxZ5Y1djzUcN1lKuNHJpUbKYS2AKRj0AjDe6mC2TI6x85z0SvQO7abdPEqZTC
MNgoeRyWrfsXfwPte2PPFUxnpn9iqyAsMi99ZAshO6S68dZI+0DJAjd13NQwXSw+cpI8IlALXQVP
NADKfU2nUvuNu9SZ9dThEM/OdEzc8uMEq15l4/p7VmPJJXww9c65zLSR8jFHkAXpoXtra3zisth7
bQcGnhw93oAkHE0W9M/76AHLdLz/+uv9Ev4HlLMmSNo3tYw8pV4Ji4ROqTnOkcpy1Lo6iYNeiYHV
NKdYg+heFGAwpn3n2Ml469tRDuy21scCrTiC5NpCqxoW+guCw4ZZXamQ1bB8VkQ8qZk70DUCmh4q
4JqtH5E3YnO7b1jK6HFbu1uiJ+UeTWBuTduHM/xItiIfMDyeDyNlWbj8bZiqK2qAQ9P9PLceHuXk
XgxgsXuYop8zPHybe/8E7upWg7yC8jDVtNoZU/yaebFoHdaVO+5oU0bWZIG19HjO/LyM42FUp+sE
f3yoMZeBIxN5ujiqmmHm39bV078TJ3yACFjbmiSdJMumWKSPmyKc1ID1zyIeZJkJOX4DbiUZb+jX
OPJLwTGczT1yhdgmoPKQi53LYgCuXzKKuV37OyJQRCxMs/itK5TU8zGs/a+xwUBZRk9k8vFE8aXY
Wd6pQmuuxFTURQ97GdM5j80B32A1uIcj8R+smLEC81GidnbLr9FX44Om2BYYX7qTibAxUedqQAHX
c0LbZ2XzvbShUdlAgMcj8B/e8qtLS37wmt5E834lWPWEzxz3/Cvhx9DZYYw+WNNz9hpLMqxkyBI4
8Snr0qBdZIsGOg/oufprx8VzCYULuZcFLW05Y9F9P2ORb6L1bxlCXQ5J89M0lc3lecALkPkfm7tj
9p8kWSQyjzQ/xC7MGUxAY7MsnYrLuQlMwWoP5Lj1tqqKazzu/Qkeg3ZPyFvqOjsT8m5oaUygzRmn
vHY9twZVMjQUWQPq+z+kmbG6itpeVyeE2ikhQaRFRyfzeQPTd5GDxs8SVKOiam8napCAIxqvPuBF
KhpUeitZoMFIlwIGxs3m9G0SWFgMSqjFsB3bWZgqKqy2gokeq+mELMB7y0KJcD4jzBiFy1fC1+PM
P9cMKhk73UJ3Re05grfdVIGyhCIlnhpG//SXKL6hyxjLr5qnpPaav0bszedjFJL2IjGU+sHH0y7k
vi5ypWVPgJOOvisSdeSQvu1P87kC4UuW2FrU/MKPC7nIa9ZFgscZ54txvBcvDHxN6YBHeAzbaZAp
QdTURhWQ7vKI6l6I4eBzW9Jfx1U9eD4yQFSqe90xzsrxS8w+TN3uzHsqpXul+qqPcnwnyqSOCfy8
H7tytsKBwJCiHHpTRHzraK/KGzOO7vDE8lCW07pIOIR2KTklCaUyOlpNjM5caBaAQHOMwxMQH684
JLPgQloD/VgG5VGj/0pjgAc5TnXmi5A/K9jnJzzFXiiQlMEItyJtQg6np4kjSYKerjU3mh7G/K/M
TR3eJ49dQomFUS0hiV30QiMloDI/vrEbliFKUmdwQEveqWlMImmH2YjIQGzXzgnlvErm8Q2uNKg0
GcCT8BQ9w3LN60hTIYL3Tcr7l3GH1hNCfk+L6MMRiyNC28B6Kq5Y07qI0lGsxRPZGjjmJJXzsTTC
ceZdNPieVKO38NFguwbvBB599z01gT4TdEqqgL/t6lyAu2yQxdOHaTOy/jpy0ba/vGOkyeimgMSr
TIUEwTQUjjCqz6Gzsh13ZF3XGrbsXEDnXCy1i59UqsTCD7nO/0E1JOIBUNOEtG99k/s3bTcJz42X
BRUrQ1S9Mqqpds50RXhsNgOmkItaRox8/IaKhkC2zFn9Y66lNo42jaMGLDUecCKAe91NOmSNlOKw
fYLJJl1FG7NrCmdgMF4lWFyOSOmNWIb+wBbQLkK8RyGFx9G0GsHhAIZhj5/3AO7kJ4A+AL3aBDWf
xFose1JqVcI+9M53VV0Pj3d5AYPvzW+q0IKrg5xLV/rbmagB2IKg0Xcu8HSKlxJNoO49GePqwK+6
ZZJSyfbhKdOQPXKtjVcJlbHnCtgLF2YutzAbeoftskrjKzS5WBLwpepHPMCDP6L8jQXlRhPTjZTk
1DXVSLOD7tAtR1zB4MUJ2WpslTJaUYt9j31luIXSsZTQ5mOMMFis265OkyvApIZcxbXSScyeWfn0
BYp2Ru9lDObNv0PXGSLhFMrPaW8NoxoViv0WAD/jxVmeQD0hBYoyAO/PQX1ZthpX0BqNiH0/AUnu
l25FfJmJeuyQLx32GAOvSomal6zgrGKZO9FK6+twSr9JYIkkXfYh/S68Pg6xYf0dysAu6TfaWQ6A
v35YetjS2xnfSHFWLjD6B1bFpDB5mymmhjOXOGQjPfB+EC8U8HZ8uCyedElEhzwLefqt4bKD2se7
y/pPJKSRFOCJ3MZI0uT8OR7gSxiMiy5nr/63bnXhmTGSjqEWcQFC3bGDcXqG6k3AojQQqm8ohEwU
Bjp5KFeBGmalBFZb1oebDQYqXv3iiwmVSZZg0+uKb+KdZX4FgASk/qzAGZ8W96Fk5fZve5GLz3lu
8aJNWRBXutgun8kzRWq/vaxd/m6+Gu2SlQWZsLKbnQdkbIcJoZVeIachFKSrSgR4qjm3HTlybCfw
O8+YPPLk+sZY7mWw1HWnibAyK6L4P7yP4XZ/HQ50iZhWQtRH/pGSDFBZROx1uGBPxxwyzkJttncI
7ONuatLcVOulx6D5hoXdiwBZsxY+ysJeCWOQm80POc2s9741NOL7TbKZYsCuTt5BIVwGqZtZJ4CH
z7ianQF2JIO/rwcHNLUI/8AEXkKSNS3bQOvoRagC/ZaaBtshPluR4BL4m5nLu4zfFel1CDFGkflv
VYIiycN3KZyQaLjKH1sV7K8XsDOgimJY4ECQNXPUVzfOQ1FBIvFvhPatMffupmG7ejKza4k9INuO
nXKLnIW1AGPXmiZla/rQj5yuQPakWf1gNXbtqzWHy9OBmZp53IIITwU5X8uegY0QhbtPmNyzWmBa
mcOoz7NfFHpU0Njr1Z05VmaQHCdWKx3Noy0BWfJceARyjNgmVxG85Vk/NnGiGPf7cdiPWNMwpuSL
ynajLq2eSkfzNW/17fcnb64kFmjuMCdwitYNT4FdWZdPoRujS70aAzUpIM9yLlzRdhNsATVdi3SP
rcsF2mRZ5VirnzGC3F9Xhydxp96rJbAQi+Dj2CVmSyuY/Nau/IxCjrXNdUTHpgofSTSXrERXCmFj
xXcunTJtWDo2KGRDvvAEfZmwKAysKJZfpb7RLxCokh2HuAmij6Z8N2RjI0bFHOGBDpuVfyBtWlh7
L9s38e1ppbdG0OQTG1oZDzD/sPhTkoUBEqW1TDwVHLiOIpQn1WUy6AdiwjFzv/HphQdb10FtinZY
u9jpoZdQ2RBSqGiRbR+6bkgiLK4jAkEjp5KEs9AP9AmB5C1OfKPG48+aFdNmD8KMAOA104+KKh8e
bbv10uyvW0ctH3lKVLBFztMYzVBdwx4JpFH67MhGn3DJeCMfZFzps4ScxJ+rhHLeq3ksMdOR9qzz
hxIKNnxwGg0BG6hfievYYJ4TboL14KByGI5W5WwpV21AiNKKcxhCzG6sBI5lsI5UqP4NMzTPBshI
JekVFTcXhs0c58eIOdh+VYFAcca3uR0mGnd7jxHoSiS01ow0sCid4VjlrbBa8/ORAlHhRpsbD2ot
n6/ZbPf79qQCB6XESfkku0l3LLIEhM9ryhW4toWy9K0Qm4Rnt9/1wDRpDxGsdxDMUsQTcGx1vEC4
myGWaEh5MjzxKlvfsS5ZVyuKc2BN67FiEuRiq6J/U2QK1/P8tbkzJ3Z8Ly8fOcU5lSlIGorNZ6uc
K7wSJ56zoHzndNd53ge4mgwwa8YSja8y9QImif2aavSKk1PUT6UFWN3troquFQ+pqZhLjPzKPjZo
RpdT8lqiAgiLU2+ClOduCmMLaYEWEHMlOh1rCZflStvFY/wx66nd8Lleds+Poo2DhTtTWJ+iOQ1s
49XCXJ9sp5Ck5EwgWzZHuDXdfyWzTvT8LVVJjvwNgegcfpuM9qj8rGB8z4JleQwdxRa2AJYoViLD
z57zFZFzSXUQy/HtKRMT0U7Jj9DzQOxtCVhZR/v0f4y7TiB/q+O7hQ2XcD1XWZ4saOU5RoKD5j8X
jFh0ED/KqBKv42S0NcwQTiHomgJhusZvYXhcIKZNaZUAV3KaKLXUdrCGf+zGIO5yXX9wd1ZD4uIq
YpJVIEkUjOR2XJ6nlxwbvV2iilYnNst23Omt1mtnrBSgjkaM/gJRggrJNdxqRk+PTDOEU6CA2syk
KPFCocCKFUGfmbE53JqTtwgW3XLLTPS8alvgMiawQ2nqWfi8ZGTLVcsghDDfS+PcsDlWrCI9jSj2
wuIOgoPOLJ1gxRh3nraUdy28FgHBJ7IR0H5kaqGX69wztM4Ii9VJ9WvUpFqqjzGyajoOUjmdhmrZ
23rXNpOAEwyxEhYCKEKhCTFbxGyNJix3ayeLxNzwB7urn5FtsIuHhj1DKmsL0iq1tcx9e/iu9Xs0
fYSzC4zP82kGRDef5HBuH/pLV8Oi+Yt+eC8mbGG1NzZR+7JvsHdPXzPPOZWjTeHnK8onW9WzTE80
B1EzLuDDPIpxa0O02SJP0Pr08HMcEIQKM6fRHOhWOuEaIJx5NmnCcII8uFMhs9vxcIMZ89Ybt7sA
9bN9nOjns5Znid6VQO2ZMrLvF8pOZrpllJfuJprdklA2ShrYfIrOB2d8L+BJEX5a9OBkZrJPtc+p
dduL/QMo2jtwjA+L897q48w/OU45Q2GAvJkhmOmjvsq5WzCcJNeq71hKAT9TpjYExkf94qRhI63c
Yve9Kx5a2J6+CzDQAmCvH2UrEGSq3A8qE4a/TN7t1WdH23YYri/jewE7M25ieEHzgQQH+4g+JgDO
YntOs81scV2b3gBe1yIwnY5SoMSpOWaG/RIVBcB0gw24Y3cPR3KQ/DOgjvNDAIwjRwR+tG24zQ0W
4xKBKzg03ztCO8mgZcGhm/1GFreazwWGhJ7btfHel+EONc/pVcNXgh18OyWaUeRYY6IDW+pff0ib
hokAbz9+GQO8JG+C9W314+JWViy6F8yTgrNw0Zw6Lv8T1L76U5AHcUmirOb4u7H5Ec4Rzm4bxeSt
YKT81GEKRTqErPAxq2DHhk0t2P5jH8evWHvwBqFlidUl7fYts3k40wKNSubqWz7l4GxLaGTdWOme
kuBGPc4KY+/bOIxSj1BMC+PdQfJTNcfY24QZTSzwwVJUGGB6RSfIxLzgE3vpT2UTtGMaUfX5qFFy
vqySXRRdWdgVo2vL+34yObioSgZhZCUOr16PiLh1EWUJLdoteamtYZMe6YMO4GOlajzcbulyaLwJ
YiC1Mhd7wvAdFdaRBh0sWgap9d66fTgFAWnOKSKKj2vJBvtcp/4zzM0CNqVMrEDE+F4Bq2YRF5Sh
1MZRQVs3IIQ0SitWEBsHjDOb4bhSCsIdKLga3ZR3WA+E26lgNHZqrgpF46dMfSS00upPjh716wzA
SVtkfSGNG36lruPKw9a8hDUSFz1+m9sB1NxxSvFJ0y1+s9PRVLfQABIcUS7FN3XraC07py8FwtyP
0qMdb9A9bjXDMyqKl7ShPMbCvkxBug98yzpSW3O9ME1YbnFV/RS4gVAzTtmY0LMIq1c6nWqpT+c3
11R5eEkXM3+mIX1hyomLLYu7JHw11UyT2dmmT4vZ3ISjOVXDT3P3iP3f4edTAckkHJDgzpcPHBRx
qpdiWf9QA53SvjB+L6TOIB0EBh6amPCowNsdxRqh2j2Gl//nBUqHY73utfIjxDQKApglVuaioozq
mV1MTe3KbMVjMsZqakAEz/LR2mSheWct0lAHXj/a3CCy98pMoV4PLpco0DuqjJBbfY8H76r/jFjq
zeznik0JlHzXzewKkPRWIwTOCdIEGElwwg8WQK2dJh+nDrK+EF1x9wD9LcXsoS3PquoyddVLiAU4
DCF3LaqojEqDkkeLC+GaM5GU52BQLq3evynQGw3syu+hFWk21wu4gDfRnDlW4y1LBIaZa2x6kUKZ
yiSgGUI7nfHP9xZ0J5Mea173Ocehdw/O2vGJIhuSQzNHUIEzozEM8VuGjatEZ9hkP04WbkKpfKeb
MqMfMbbpJPfLHRKZO1J0Irkn60llO8akxAHCSe7RwKsxZPZ0n/hlhBfY9rAFJ4EmaBzff4QOfzB/
mLTpagsvkoUodZXOJfl+r9GKC19m7OhrndVMLzQ4vVg0m8mN8oLLlZgYjd9i3ZzaS0PuCD3ciE1p
tqCFrdZnx7VXRLauFgcmCTD/cmXe5cSKVSP3s4iOITPfsqsci6tae8nhekMp7wWlg++Xok+vKmJP
VhZoqODgg7VOvjDKR4rmqKYwy2KO02jQaZhjFXexaykQPdLFJ2hkobV0ntvl2LNFv9tOVQ2JLG4/
qBUoNhsejlizNn+6vbfhFR16g7nogghpGKs+aC2b+gly0VYno++0LMDa8IByfhQkV/KWD5V2dO1m
eFbBD1JWzdvQJcwx6PTkH0M+ipXyr7ne8w7kgfSwDlLdJK8Ngraeaii4l2qVKV749eJgXA/Gy7AA
YCDrqEa256olJ/g+BWmPWHslbMyxSUHpAah9OuSXIZO9m9YeRINHkpxc7anRwRB3b+wn9XtdBwfG
4YOr0YAd7D+uluxmKQHxavlpxFnhv3emzfOo9TI+g2Qm/h421IYGQ+bnjd1xI/+QwIpUK+5BQn24
imMRXlST2kQKmn+loge/89TG2dTtlbslaoaCHntCqt4e5QkNA4n0RrlklneVDrbvafgX0HNSTXPA
vBE/6f1sGDTcR37WDbGef84M2b4G3PsaYX0Ys+epiprG6ILnWugRRU6Ymhyu2A4XZECgYL7bkUs/
83Dgysm2PcmrCgcV8A/+kyhtriUr8fcXY4MMMVUxovhrTV+KcEGkd9X6LvuDVTq9SfSqmci09AbX
wcJy1uBLPoBWfRoAGn+hqx5n52NlnFMHMjX3F+jjUgUPdcWHbp3Z+nrLd63CsEEb4UD+b4NswR+y
3jP3BV84m+nk++XFOtlyV8D87/w4dNrWNYZKjs49d+YuMIHCSjHbRDzsWsnHjACEy5g/oiZMCwlj
BuzUOQTnKQom9ud0ob2Z8zkaUrSZdbCnPuA5iA8Oiyl1I8nigBQK50dLBy4XiImKC2GuuQKXKCnt
atSuks6dBkzNMbS/U2OvaTN8dDLShTglmR98WNRcj+GjcriJ7p+/ODlCpDR6StzP6AF7B1zI/VCk
ZP+ynOuA2JFMqRhwQNPn3/vMUrFKpMr3QCzz/RAb9fbXG66bG6bODriFoP5P5NUlHEIM/3nPOfbi
pb0vH5FaIrnDKmwhA1yb1hPaN+G4UdDDgqkNhTROgCV2yw5BIlHenbhGrLL5c7qyfhYHMwWsr0jv
kN0gQz3xlqwNPTTtjlEAUVCyzdCVWHNN6GDAfqNlRaMBFOAVCykBhfso9mFr2oM4dLiXXOAOaGuW
7ZlDRZQDpJrbCNyCLl8VgcXRIvamTGTV+AlhcBhSqf/jeulsZCZvh+H9Aajw5iwAuqbA4fcHo3xe
zEXbMAl37ZT511QTItPJt6KS5jJ5IDa2xyuX+aFn+DpTShHjOUFld1nzM72wA66XlPEWZC1Pv3lJ
ri3AE5jLe1Z4ssb87AIeBxJ8wGSVLYwheLT2KRBMvj26+6XACsrO6L4l3CSJbfZI263eUJGfADEx
Mn9gDtr2zumhYMLGQIVUBst71iIhbY6rJY5yUlIoayx0jLv9xZFeLNklOmJn/6LWW9nANGtXRX+U
ckEz09DXDxuoGM0qMIQlKnm/iPodPLl2SNO41uXGyZzpm8fSDVvkjkugyEgNStr6U9mtz8mbcdOa
sw95xOpLI4NyLZSCxNqVn7SUY+yd5zhcdkYbH4uZrATtz2aF68uxR6kn7Mu4GHHTY9Q8wv+XZNPl
JVLKv7MW5ggOtnsUG6/576RjnpbdruvohmkTbLifxL/mdmmtuVHbS2KiO1ASkIUw0NAX3oNopZLY
IcOOyb7Dc+Me4BZ64uYuSI5q+dcphG7I6yRRglcxS6YsdEE3Y/dc80MIpP4AapKtab8uL/FOSnas
RnIowVTNs7QtfTh5GQpIbm5G9kAi9nvdlQB9JF8BSUNy0hcJdC4hFHgY5xE1AG6mwG0oN7Q9S619
igIVfY+GGHexgaSOQgK0vQhvuDZosgP6+dQzdDxRho/nrIBym/HO1GejHQj7RTBrQGO1HvtHzZEh
TyY3rPD9NercN1otaBganUwFUuNwsMc3BDjtEfS2NmJclj1tAgEVDL41gNGxyInWCLRcaRqUhrxk
F0udyM3AyMf109MUsgexsoWk+VnDQTk6WSX/WVHdzblKcQUJjWYetxKyBQvtVoNl81l32X2O4oWb
XcXM675ujIoser1wSIwXpVG89ur1bDnQxHob8vsf6lR+bojwlhBAuJrdJ6s4Ws+HFp33bula5JuH
rQy9MVAXQduKyNiKVbNBNaRX7/b3ITMV/6F6LfrSvLRw2Fd2UdpgpM8/KT2ugtjgaJGYiCFR8uBT
bRk+TUoJ2AMCOmAs5FhFh1JYAF67WY01nJLvvzl8sQ5wF8AvRWZwgWXP8KgNie5+2eHqNZXYi9QT
+tHaWmW70jqLOyvkumet2adeMIHgBSxdY4tk5oF0MxENmhpCezigbMVgVet0+jObhvvQR71t2Z7j
/667bHJpQvKfkZ7gG812XQz84q98x1VzFDPIxDYGvF5Berwgp+0HQD4D7EtOpPzHVo3YDz9lCdg8
+ovUlZcb8XQGMwlXy6UNhRJFr5Y70M5CmodbCKNGSReQSPjjZUoLw9c1RmAdcLGrPXFl0WC631IH
gKPNifyW+qqj1vhk4amyrmO+CgBA5mDOpaCSti29zF7mW5lSARVjV6Xxf9mKB/e0Wh3qzV0t/JYI
4cVuKLhVmE5SKvtYTG02XlDN0SltPEo4WwDTCED0Ov8eFRTFGY/5zMtMYTf0mhAI3l8YAiE0pU7M
h/pSGf0im9h6FObyVlM5fMySbn7eG5kOpr1XT3v5Coabvl34um79DYIdCAyUuNlLuNi/aWJQYp1w
8FrNuFJbnhMGDypU2b9ljMMV/9IhCagl/Dm8B3LGehUaT5BJDY4CI8I1uHCDiJXBNqJGrQeuCCJn
DOej7ojGTBdqDf3H7mrRPYAZoIJBIl9zTgrDgfSjXmMVExoVSVIZBE/57tY+/f51hdJaVAXsv6eM
aRHNukQDZbXW0dUM7F/bda6Frx7RvfNnkSIUtFP5AkXOaSe+YUQbvBsT8HLX9bO4WXRMMRpkNQ/L
QpnYDyBGsRImRXDrBwvYlymaDid4EyaboA5pDB0etRUvz0b+m1/GSEg9Nl2MN7nSLNwvwasgA7/0
wB+82ejBe1BrfTiLLcdbkq9fHcmbHrl75PYUlwYUbLHve3zehsC4JRWNNJZNlrO/94d19ZNEauQe
hfZ6kdXdcHVc2tu5radWRtvooki/NvZBkxohanPKGZKDp7djxwzeI+eFAaRPakD71xLupepekpOA
Fs0LFB7BVqX4SOVdKke0W0ScAi8gcYsgdbcOJi8BWw/ZP6jR123aTGWN7aZ5PkrRBELinSaxhDmN
TEsJJJ2yYsh4dZtj7FGPgRE7tt3bZ6E0YOC/YmzfgFIl2582eWoml2VJOCGmxXtN9vd9lvzzQCsC
tFlE0WZwdxJrPW6JECN/k46CeI4P29hYnNNnkvVSSSQ1dUudrlNpkSIyknUxpqycibxqFiI0GsC/
OSUUIuBwjaXf/rioaotPqA3rhOkAOl7LqQJzwNeUd0UIIoNnxJiRWuV4ZF8Lm8hkAGuLFzsvQrlU
pOb7W1Ndosnq6DQI41RmLxKVhkENjTp8zFVn1ShuDoVxBjVA83VrsGTxOLb1pxPUer3YvpP8/AFw
xDkBFK0Ns5zmc+yHpmfC7Yo9Q6lwBm1VWEsokfZSH6m+UqndDVE7tyYPKiJZ7uXwlEloMT1+jVEL
ozru6mEIr8lh6ePnmrhR9mD8fJgLzSsAcy4OyLY/CJZM1UauyHyMimN8CgC5PKXuOK2JeYiSHSBU
dWrGJv1e0hURbl+/FWvd1pRZea/2HqVRasmx9hR2YNpbXpffMvwrBfJpWauzgzmUmHTDD6Bk7ALg
ov5jqGT5dC6mUXlVw18tp3EyXQW45RrKFdCflb1YXGhGuNKsJwS8sSNUWFooEgybbFzx9+5HmKPf
XS4cxgrEaZADRspja/2hE7OEEEGusYxUwU7dWUkwXxyHrz0bt5IO8sHXTOtfmUs3HkIET28bExi9
a5O9QQKXE77GnOhVSVW5r6ylgjsrWeR6JbW5iGkuc16tReKr3Gl1Iiy+j337eqoZ38/AwZYx0AN6
xJk3JSvOB0x07fqmVNK8cf6xzspWaVqc97YvA1MqvIJNEcoOQr2zAPKKYLb4J791yZuaViG0IO5/
9SVkw8Cw+M4NA57D5gApacTZ7E2xXj53Ui98w366abGfReTdSIYp3i4njfB7r2E3bSOzLhTHs3Xa
3iDkAD3hl8LtZCsf5z1hb1WwZwIjWHOf5qJ6RW3l8wOR3oh2/+KCrmzJhrNiHqlEGXAJH+edyk95
UaYVC+QF7o/9Svx1MAYuGD9o6p3AflYannPzqqmJDAy2tx1TYcbccl0zZG4cu9/uBTo2+x/yR8sT
BA3A9ZqbdDXQVyAEG+uFwhHUR/v25HG17cGJASeT5GcCZFBvYqb1f2mofLm7klg2JQ4iHnBSWoSs
NlP37SeIGSfluEB0cmoTxWgvhWldBjj/qhGO4wfkLvQ6jPtg3vfuw3LYIPxMFQqJ4n35n6lio2WZ
35/QXjFrl83fbPUgiJMgmv7aX4F+gy2ApKLkLv0rfLSxfRFalKJ6c+obZgvJiis0JEWy+Nt+pxH+
5mKgcr1Nk3I2VNaVvcj21l7n1EYiNUH57L24ZPaYyhvOqQ61W1T2y4AOgVH+yIvvV8yQ7RyKLhnY
9wd31wGmBoGh28WMcEitjLkot9hwIIQwjH3aL0GHW9sPMq36V7j6FEzjgQZoOI7mNFeYBbp2rMkd
9raq/qoFQcVhTS/54jp5dp75//IZyHcaOguULCGCZGAuAVBYcbC7kaVQM1aeLUPvid/zPwu/nuAu
NloHUtT/Zdg4NRqrxrXZI8MrEcA5ttqaDAGFlqvtgiWOFXtuxLZ7qvoaVUtQhUOuxkNuQJkOBOsd
zKqzDJu+371IWlNpKXUtQTyWIVirReWbOpwowFtoMihNZiSwEcmoUr6CUpulRpD2JcWcPJ2O7UVt
GSLJD04c0EVba0AsYoAqh2sEKg7XyiBgCfZXeHeEvXu94nXVtuia8bRpmGuefzX9xARBOmjGMHOh
/iAfLZ2Qft1t6557GNhjFfj/3FxS0OogWj1LIa3lMnBzvAVSq2aO01khXVosDNBjE+E9iU91IInH
5UwBF5mp/c+yNJ+T2hAlGBb4px8FCJoiILNVfkkzTOPKJbfHq2v11QBfqHcXIO3Zuw0JL4cNJCei
N72F9PK4M5daveTUaJTpAif5IzRjuarZtHBPbZjz1MBiFTxh+SQ/L6HKMmC5mMjYPfSC3Dpieb95
fQly8AAuPZjq/9nVyaWv9vDqT7Con5Hl4DzOxNRbXfoiV2LaLon619cK52HG8TWPkNTHHQd5mqSl
BkdrzBw9e8lMXO477JIwCR2FwrPby9CNJn8MKv0GG3VgEh4ssrF27aDQfjPkX/Jf0jF8nDrs5ETv
NLAGxP7UpC7B7aGZSBgD0sjha7v76qfKzlOwc7LqZxcTOBco/joOwQj6XA6a3nr0IW9QIoxsvVdw
GmTM5Ccis43n1InOVS2ZQOVO8Mu/7Sgqs6I5OLEZTrMrRLOYgcYB0vLNKZlGIXMXL8H/5GOBMPKS
UJSXkpnXIYFf4YadJ2EgSR3mRW2Sd3/AQdeKz4WcXtu8d9deu6SYzIf+foqVe+DXzsRk4erC7n2Y
iv5+WEUKuWKGL2OfIl4N7NUhxf3bQA9Hwn5Q3blsHI/WVlPtxaJkPnlxO8SRDSLKarLuM+bN5ySi
Yllwtp+b5lWRN7sOdpMQm44sGdgkTE7+akg3AubNgVnJQgzb69dfUu/Tg2314OT6bfI3q2/pGahR
7YKrSjeXu4QjwdyPRLDKBPCBzjgnNtrOCWzKekVAbaeNw+bdKGCnIxIa+5++CcIQHJyh61fgvwLj
5tBezwdAONjKCanA+mH5EpoaVzMGyMzS6h8BwoitxWbafA12a85IUTYSrA8OPDDetSUm2PD4kSN1
c+i4G3vmjlqEbBrHu71EnxoegLFqAyqxHEvc/jKziGrQkrna2IESUeqNZWHMWcwdQ67Nj9XW6l0p
jvl8PiGlAHj2fMtu38GQPwrXRbDRTXJ6holI5YnI+fTISpk8MMEoYLPLa1zXGSQx2bGn2PRLDanZ
rZnfzUXqhjvna5P6zAFcesHa6ytFFe8kMmukBJwLrQ3JNfI1W5KaMZaRJXyzyZeHDsdsxyEPzDUX
JVWqz7uB9XMwL5/YNxrzyzxAkg+V2FQNFTxNB3HiJh2s3UMzZfbW82cACPrX8MLDU0XOZsSTGOg/
N+KFTDZzodIB1vAFJGT3S7AYviEn6KtXb2/eF1XWr76vkd7N4BODMVoRf9J5gpxASNbLDhKXpzW9
WWn5xjmMZT/wOXoKM4gBC1fj3ZyC6W+s6V0P6TuCLr0selt7vws3FySg2AJBh9lhUlZb0C5j7SWT
iFvt/QftSBMdM9ULHgXoQ91cuM/MuaTi0aqQKBtQ3Rmzw25qCQVy5/4rl6JYBmIjrtO3MhTdxo3e
7itMyDGDg4Q4xGqhuovZeUkInvsx6hD7D5bwwZnqsljo/xIdFqbvvrB599Adn4Yp/LGLBjWc7IJo
Vprrz4tdkimY77FL93lsS/1ClP5Teq/33ERXA9vI64bDJSp9lHiacY0XKGpqZZ3C5ckqn+Acfik0
dfkhGM+vhh8SONxDWX2w+ck0T9SUjJWryJUNYLVSCVtxzCuaAaCBqt2Yst72SAq9evMgxskMYJB/
agreCZTU84jMsXK+5s2I4y31Jz+M7VA8TG+QjvYEkYerD3W/VB+vnaBxI04Bn0F/9IvFxjZg3Ivv
1IrdSQvDgsZnMX5dayYAlKAH1IXhHbAahjB3GyKIeeZz4H7Li7MOfn798TJ4zIUTCp8xFqnxJAbs
DmqYX5/B4/IwPbr9A4dzWSZRU2F5Y2nUCDH/BDHPUd1eA7uewmsiYSgUmH1EoNNLgY6Gvy9TIOhh
8p+oTcInRci1izLQnH5GSTj7ixssuO9puNRJjHBCDBABUt75xlpTbYbWbCTApS267s1KAEJf5f9o
4hbcot1HUYyKuhlBOU1yv5wBKhV0sMJnAHw/IzzNgNNmVy0+6WXsej21rXX+riHGnr3nV/JDa5OY
fYpwEvRw/uytEyeJclyiDxE3i08WSjNfRPawysR8sd/VNgB7e8YnC54JWZ4uld2savWvoyM7FhS4
DjG/rC8nY1/Zw4//qlg0eZpPi/wDkTkQLxV05DijI6fpYMGCg5hBmusrp2Urj2OkY0pgIx5zTxKS
HPK5ybmcRlbWxQVPghUojUaBL7YNb0jZ9jLQv+TfhtsELwargZCu3h37zhzAIAVPrSWGpOtEF87C
djupeZmHeGRF0Scot9kSwl4jWaZGVOioDgBm1CEa8reDiWJms7JStNfF7QjRmC8bEKnO2olRgJkS
7rdSEsFzy1KjImbxASl+mkonOa8N/i9Jqqm44WkTebEYtb4FrVgJcWjyat4xLRLCQCjk9XXsQyMY
HH94y8M68kAf1210ECOWT0smPTTuyttCAwGmz+lBrkLni/Xgpi2NJGQD1SbawDWzXyFakBaOyXZJ
vF6f4khkDg8oDWcIF5EKUptBhhvphuyrUGiRcG1UeKaoC+KVT1pRyE5+bkNoMVMMtMcTz3sQXQxZ
4cw3VU3Xw2cjb+RU70rwibVR4DsT9at4XTNwgPxU0ZHOTvI2NnmpIkeECRD8N03O5FaD81GOQdhR
twcOMlbOt386HmDblfcqAiJ6c5BDyZ9/AiHfvtxsHqHhJ4+dTywKlocq+oyT2wV2zxxskAM34UI5
QO6iE9L3a6QmZBJ9loe0MjQx+KKuIENUpm3so2bMCwhE9cmZ+YdAbU2SCm2nJRR89ys3FvPZU7ey
Yo/wZ8/TpAcZOWb9yx0crPuOmbx4pYZedT7z+ZU9t35I5E2t3QaZXkuDK5MHM5vjO9Ze/n3knYbq
+XmWIkLCrFqCOXPhiC4UUhMty0Usgfn3DiGDjzcRKrzW71AiPb0SckOLYFDBsmsk6bHfx/nQ87WK
SYOIB65zY9rMIpgddixyZhgLJMiVDaNRp6BuOITK3nhi7yL4KIUvrhhArZWhpu3aVzZcS5DmaF2t
p85Drw+azAF6m0S/V6c+Nzc6qcP8riDdRqk5bf94sh07b8nvwdmBnkdUUnx7q7ibbM36dWWAZNwY
4TbdVVEFw0iXfLjcNQG+ATjjstc+h84ww0BOKYXMld8oyH3W5kEUKgm0VruGsQZwdK/kk5ZamtL9
v6CKw04IbeatrbqbJKcnuxcgYIl0x8IZXnRRIb4YuoPQkP4u3uyXtrRCPTRUU1WM9eJC4nIhFdYN
NgN4zkaN6go4j13FOcVAr4hNoZIu9Sef0VJgZk5mkEOfVYSYQ5C3DNk4s1wh93kR+By5RjnPcNK1
/Sztt0k0CNK7uKXIcQlTmPQVB2C4hxQEjnZxXsedXcayLmLZfZDP31sw0FzzrM0XSMJw0yoFRUT5
OGxtkUIs+RMZ5EEGvvvcwqg8zxzwuu2q8P9gPyt7+R3Cuv3qVoliSiE3SpIixhdbJVcJ4zV2bubj
SZz64wYXodVn9eMJ4+ewxvQ0UOJoqct/e4C6dbu6upU/QeVxjVVv0mA4200D/5VFn/CZz3vj1eS5
0bP3P4mvvx+20IJHe80MXaqMOxqF0cV/wzmszRgcsqyYk4aWsG1LAQps3sxgPJV84rwr3UsJrzSt
yZFDY32ki8+LeMdzZSNceIgUqRBEkDLjZeDQ6FNfTRMDRbYw/fi9YlMRNk6eZv+Tyv8FTYXdXASM
gaXRJK49OPVOxTNxuqHRMZI0EuLB5wRP9suxA4Gr1xzwjX/QgjZ0HSSg+0nHGdfP5BrVuv0eLUvd
u+JiJYTIrzrJuof3pq2Mu+MhZI6Ur54PYwsHIx+nyEsOFskD2nGc6FnCvsysMo7GyC4BpKpPVCFQ
+zcpnaGSNw41fspLQ4sCNfY2D4VY7lI2Yyu+jxBvAmlc1dh/Ap+emj4oY6jhYf0Y5F7Z9N/htIJy
9+rKLEY/ACHNjDz2FYZopBHZd0ORftm3c6Gzn5cUJErbndzK6gqaB0uJogt9hsrqc/jpeRpIF6vN
Rksiv5D8x+2YGj0omYhTZki6rESKLg8AQIlNeaLASfC1XxN764iUkElgD6sM6TCMx6QllnlAP3yJ
EaqkpG9rPJ0fBud+dd/lkMIBW6dKo6LMH6WWJbS63UhqQ0DuJZPfQLwaFzsZnmQ6Iu5WRVesbtOh
eMljTuvnhiklpCAw3aDf91t0ixgxwcnEEHdgEnDDWMMIweXgwD8VyqemueAbTKbo6v4yKtlxll9e
m+8yjc0RT7ILXFj1UjvjFJs8wbJWUf5KY26ZmMFKWaYlLEwMbFM4LDajxSRHiMRZiFxZhWeWv/Az
8v8JKJX07K9yl3MZ+yr9D4U4rX5YkXSiadVgR4e73VUWK8k+XtLp1LO969TgL83xn8RKFMCpHCc6
///59A3c77HXexyhiNpjL69aQH8m5T+ojVKCj/to5Oq2pUZS21fTpAEDmB/N3YMXB8ATwu+NwUqm
BW+9BZA8RmDz7qUZFIvE2rxiJP1Q1U75CO96bL9c72rLjZQIN59cm4SHpRxJDoE/fqNvXx+0etDz
Rx6kkTXy3AbITTbVSPvlRgnyrR1tHX/R6R3qwE2Y4zPlsL2l+SuDkIEZB8YXq24NDXzEqRQbpR7U
FChm7QvSgVqQ5KMUnw6PsjE44rzt9t9jBGQS51i89e/n8JdouzNOny4LnaHSACC3DkRUhxA546tH
X3j8ysRTI77TnhgckOyb5w822/A1fU4vlv1YAqNnm/w7rp1nbbCxorn/CjS/a3SyT4FqxDaz00P9
tOQVGMKmknjauE0xN9K/UNRP4ARd4wdEOkm0MrFJqueZtGLBoVkjFFbswlF7VmHyeW86tPGJ3F5h
Knhv9Lte8eCUJhH0ZFnvTni6xEO2u5v6KgffnVNd/qYeDShivZRmINHzCO2HNBnOS2AIQC7qL8wQ
iwXAk+BsQgoQAFtjMMuhAAbVgQ5P/s/RNqlSi3ufCJ1H37ADFIxtf8pPJ4fJSCcwiUEAFaBAme3L
mr+YJkoE563W0P4z84NOIkgpkd6Td1MzZTq7VJY4Elpne6dYcyBjko5YeYs41YuLHwo6IfzAiKT7
vzSjJr5l5EgtvEbeMDeoPU3DILOOsdTKxxDQmbmbFc8Zjd30yAt1YjtEqThQj+dt8UW0IXXM23+B
ApSjfF4QFFg+nAR3CkJ2U3rWeX7/WEgBeGLN5TLoDPU07AqjWWLovYiqksXJM0ynE5Gc916V5f3V
TLflXOOJZ1tp4Mt6WuyqpAwRHVfozlQtFVqOWK3R7xNQrFwGxzkhRpZ+74zstbzcm6N8GM/UuZyo
NIDizjEJbxg22jmDV+fkH7mM2xhMwB0BJQxYNT5Kp8D6J8v/Vsq59n9Xa25P7oyKrGiTXb+a+K7n
LHEl+BG9GtN7iwgWukR148CcZHC5sTbmQqm3kACjyIvjno7XFUgD0trt437ZNU+DtoYrvEW9B1dT
UX/9qSb0Wh99FzSdNV5a2kvz01swFUUoxcBVjLEh94qLKB8HNcysNXReEufNTtxOBqydSnEgwyTd
GmS6AfxBVQMJ3VT+yGBbrxNIHCUHpDfWVTvUx6OEPWkuppuF2eAtFEmPRt/7R48sF8tEvbO4Sw6L
StjT+YjXi2peftaQADnUTdKWHQ0ImX6hLscIVqZf4knT30STzqt5iSdzxFDuTbCS3ZEAD1lDf/t6
ydgGDepZqnIO6+OSsoehY2pN7485Vn+j4HJfSN83ywBta0qLIxCmBMR71b0p/lmxqMAw5wAjfK7A
J5XVZEjNzBbuMFC55I20uHQTajN/xCseanSdv4xXHzgPkTP99sSCoslpvk6RQEzk09+JkxMpHqLB
bkrPTvnx9TGnrihyUK7zyFkarYS/ONWJjt69uMqxzqbwNOZAtP/ktz4UMIT4akP+DnPXGHE9JoR/
fdiwfroXcxm8g9Vf8+VlWDvaJUCACRjGjajlnPP5nip0mkp03r7Y23TeR8L2rNqcCJjpUPtRGMnY
hEmGLUhirlQgRguBWwoLfcBWMYb6MdahkDD8QNOMJXARUkQ8MQlHdgropkS6gAh6sifNJ2mQEICP
EeV9NdiKZ3hEFWFxuKGNpk+Xh2lkZ1qg1f8pwhpT5rU/1TvO75YxD9eQh4bhe2es4Us14iTHzoQM
nsKLT0sEdLXv7y82zIlwBSVNdhZTL0Sdk078vk6E2GHrlcudgGg2YY6/0C7LvzPAAeNghQB21aDs
BOAg1Iuu0z8MklzzL8Lzqm6WtaXpAO+Vp6a/GSNwsjbzTIyXvBYv6wT0w2ukvz7d7cXsSyoZMeD/
LY/l0mLFtEoQT5SqNNd+HUsgAVjGWrZbDM+p7lyvaGzdMiff6+WwRNQBZJLWnrKswO8G4Kdsrbro
z8cDEO2wLfG44WUUNNkHaylnlnJgLFq6K3nzrBMt8npht6HcDLqRUz+1ZXzmc7fyavxIDjXUw61W
4B4NzVlJkgpOtX7o3jz9HbqOXTR0daIC8imzqUHrSOLWHES8QmfBRqNQ3ChFdD8/+/OVAB1e+A0p
j9PfCTDYk1O2x9IQ2qMz4vRO9pElfckUSjwh3Qd5hEdvuXJDQm02SHCeefXtu/4MG6dcURAMgmrN
eK5j186kUy1diyxMtdVxis7dh942F+F6U6taouBwD7KVgCNKgsOvXGmnfeuKNZPmGd7kvaTJzo8B
/g3ZIDpkVMO/M9gc/2CvEqNZeytbH4Ey45XGZoAtNXOirRJn3luABPrki6mwbI0rzi96qZDzoHSR
cbylu9mInlSpE1UmF7kPmOe8uN5yyZ2WPRAlmnIKn0+4Isf4JUS3pS/2qtzOxHIIJ1C/xGDHJLXk
Pabie4lpMnjZyPJUZimaoFywi3bFrsWpCDVkIdksYj1SNdbRNOI0BQVug1k75A+VP7mR9YzwbUwj
vIg7EtxstT4hBIZe55Jq9KJsGdaZ4Pgz0SRsOREQVx/Uy0oMZB0ThJgFqHdUIU/5p67FBaifFIKO
cC1UzW/j+4loYkPMp3CZsz1fKV66a7J+P5f+A9IO+tVq2lcFVVMkFNb/JcBKEKsDIpFtsVSPs8Bp
ZDtA+1pLD3t1KWixm2qcmHmezZbfExLAAs2oBP6uT4awIj8dIQnnnFi3ZJ9Vcp7D/KDR94Gjku1H
JGYdt80N7WLWWNHwFTM3s9/HKPijv0Z95p4qb21tF7OxkQNjwgu1jn72kkNyALW76MC8mGYcuS6T
ZbxcN+6kN7P6cJ7xDJZiZ7G5uziLVgsZrLbg+lLv6p6Ui878ZYLtcP/3ZzGrAs8P0drQ1Tp+PQV0
IOkd1SzQOJkMEbVdpRAlobs5W9qJ34SsdnRYJxokCkf3IWcLRPdTcpcEBVg3rigT2ltVg9RMvaAW
j9gbeiX3e1uGF4YAQtePtS1fKurcnMoTEmW4Lz6U/3eM0QTw0Z5y3mQNLjQ+2GzltvPCjKYyM1e8
lmvZ0GoaVdoB/kz0/EGiXc0iS1J+HzqvWNW3Up7a7/iImZv6cLdAZ+8rQSMtMSHo/WWs0tZgCUEP
0BMhRmOOr+r6YmRNgfkeCb1AedueaRQIXM+o4gKe3uXIBFPEp48boG/7gc/qFbycVYwwiqJOjZAh
e/oLmEvyr5o+SSD//bWYsr3qU2I/Xk2G5p1v09EP9tnOqOHPCQJCU/q+qs/YKvvQ7PXtw+wdjvZf
NGLnFvam4K17//8fgosbfAM+gJ7dAn7vypWgFDF/kTJKHaITjLlxQRUZPfkiIGg7o/lP5ifxVUzX
THPgIHyvBXevqG940jUbGEscE4ROGRAipPrA/rqB4W9tyiIwaLEPEczvkXPGs6Xz7Ys7+//CNkuy
4MT52HwghTxpDChBti1H+XQqvni8xN8LHzw2uzLbYI1ncum+5a2MEfiVHTMf7Ff24D5KslEcfljZ
vUDELThauKmdjg/Q/0tCE0ksjIzmZ7z2PSvX4j6JammfXjHR0m4RMXG8btYZu2Gt02Nes6+hmBAl
dydkRZOYBAjEn66vAV1wZlaVlm65QijgPraDyKRB8A2MkccA94eBwCGBCm4n3c4mHsd6toXx7EjZ
HXivBtODWRk1vHsMybQgcbSuFkbbHLkFOKHTtMlvEoNDSkUsSbav89Z3/PmKawZxFveC1tMt3MA2
ZdVjWvLrOYiWy6cW/iz88QiRV8uLdsc+6Fm9Nc1jCSLSKcLOVTgnD+v1KeIncMyuUQkzEKLml72v
KFMtlOn2NY9S4XJ2kCKPEzUIs05L7/AaVDx2LhMh4fgviwNouzqdcquNe8FDfyx/b6lVCF9fRI+d
V7CMCv+Gt2WAbUeU/jt7uTKiatrQYIDSv5aUwtkDHb8KO3I1cnoW6sSUGm1GnaWpq7ijtedLnGFm
EKRFey2CvBcCyQ8fO3VyGv7XcjYvobmDWb+EcGUUURKET96y7fNaPkez9ks5yOruYmPAHY7aQHka
xJziX7TBRiilCl8cHYqxLKBw4xox/6qdGYys0DmnuqdYjUFTYX0+O+UIiqhHIpS/F2yDBBLhpTIh
xN7nFLd/qBDRsB3rN21sEiTv13KHyI4TvRdtGAWdirfACiM6XJm8VcNXY4vxd9L4O3/qM7v0lMBV
nK89CZsX24hM6BdyBm+ddXJwIJWOggZyC7s/2LBdFDWcEdREpk+HR1nIHeifQimt9BcKqWXFBJ5O
fd9ou77iEmo90tlfJbs6lVh4GIT17KA0FCwZORCsukha194YI0NXwXWJ2zO8ZD8PHPVKs1tnIIw4
byEXLMzMQ2MtEmvs7HW2A+hd8HMkwo8h/YRgRCzpaShJT3dIDMYF3TasHwjcgNUBSCs4QiwVg2wK
2LQF2sZEv9dO0zz4dn01+dVWnGw1zwZtyzI0OfaFb/5s/Gik8EXrq4OZyJ61RmsuL4uyxtSWcZw3
t6dVcixV90krr3kMFg7T5R6qA3utF4U/wIIqX6X40xBvuBhiM7uARqFWtmH+1fxBTxtKOVeGzbn0
zIDStISYeWCqlwN6rxw++2iXXADiLIr4liHFXLVP5m/GfhUI7C5jFm+aSpHQAJyfSAKRKE2R+at7
heVb1BMeyIKK8xdlF1JOeEBOIXbfzw44QoPPULirxHVCDzPcRVp8SHVvSpbVHdwfEwGOzK7T1nxQ
rPWNIl+2oRrx9TdPbx/fagiIqDw3Rm7CPD27p5YPRP7xVXrbvsjFbGt1Qxbkuz1ENJRhOnhTDt2n
6Tvzfj6pkymOjdK2tsRJALRm0r/FniXAAdGeXKFK+g3l9LruICuSb7f8bjKFrMusUYO0X2xiLrzM
CB7Q0o+DPY1a2KclCRXav+IvK+WDc/sXWUMFi9KnhMgwb97RNzK8znIQUmVX78O4Wa/YjIqhBq+M
yQHh+Q40g67/9/98FlGSi2N2HD3NZd+s5h+C6wXt3Eh4xBoW+ol0wb4lKP1xs2FZJM1mIQe4zvqR
URRs+AtQdHwGe1i/lVOEmdmlrP63HKJ8dnlurWObqIiEvWpr0A/mqFMIQEjfccyMk4jy3tYY0HAu
bdP8aFcGn4b2TipUbdClOqXSRyB2nKTBsdtlJNMsDGRJhsLNXu3zJdlt5WT6JQ18dvPG5IeZX+mw
EXoJ99U4xa1rwerSj6qzxP+v5fcV74fo+id0VQmdFRG7/uq2ZUI6WBBBsp4WwsVak1zg6cl/LDNR
K+TFiIx7zxzlqvAnvO47VmOxNWi2ELAoDYJY83LGzuFz5YIR4Ra2luPrTxXubY4slyuSIUH5fIOK
V2N18I1q1nh8vBtEAGDgT6G+w+gySZ8eYHwO1dJheBW2T0NzPqspwzkff/mUyMTfT9TJjE0H3fEt
aTwWx0lWecJBFl2hu4/4eWSsNdk19KVpsXva2nGEmaNm5W8MU27b/Ff29h5BxvajUwsC3UYs9cp6
v/CDSIGBN6DrlAz3rEHJpmyt90l30xZT4Qi7DXPvX8N5NOanRt6pNu9iLxaFOxpXFL/0dZeXSkxS
r3wjZlLi/zeS7oo7octb4l0j/y6JD3U/oh3iwkTp9M2bHUQi18vtXK8DWEs9opMaU4sW54vXeyTZ
bm/WxTtc87KgnPI1j84YbOJgXDcn0pqXaS3JSJspybPKXw3O5LsNJTKR1WuocxsBNor54Sg7lA6h
Q4zWikOuqzGa+Z4lewmqYHuJ0c10ssO6+q8WIBjbbMSqttcv6DSMUuGUvHg6njCr6dnZSWfhls10
nzBmHm2cwjwZbHOm8zIiFMPQcVZcL8hv67NIr1ACn0f2sx/Jv3+htzUKglLN21IoQW4gOzRonvu2
ZCMPJ0XM5bxU94wudi0eXM1CMbK0iCN/u4JCe2V8UC/cKjUGWydqFvqlNdS/TWUe4KZslQuhUBC6
tuiD922FMqSSkudseAJC1e5O6n4Yylmqo7WXVNVQmBLZGyPC1WESH2KoPkFJ2Pr2nY80PvFgDB0n
zpJZEZZxC+9B0aL2NqAyHKgB/ko28eeP9zK3UeWfcIH4Yo1ODgWikDNvE05iQW34Afbi12m65l01
ydNciLpzKLb0S/WV7y03OmySZdh5s4F3nNLEMV4fuUf1RUokJysW2ioNz2abKEk8D6petDJnAbaD
t2Nen0+QAQ1SIRf25AEro64mvHXPP4n1DdHoPfKLvnKQcUmDXfmCWVOZb9PEfBU/HFmBHXaP0PCp
5cWlTWMAq618g+8eyVRiiXtBpoo7zjUxozhPKsnTOTNVdBd0ueJtX0pCdHcc2Z1rLRQrbTW5UH4U
0VLlVrKRz9BV8z72rDWTZnSpjzsA16u4kbL239yJTKMr65cU1YtTwCucFe1EFFPrMoqEMI5YC670
CVRgD6DZYftfWw++BqldU4gsvwW0ZC5VKHwP1H+DqRcAjT9vHdJ66uizpWK4RaERfrEIlZCAjEq+
D6L2ZFz3jssXMdzSlxkLJT2FEZjs/juY4grilVXiQvQgb4WA8QS3rsCl9IKpNHe0PETixNPdD3XA
mR0YICkK3MTkv/M51CAQD92rlMkpsEHwrrPMzSdeyU/OOkQuBpYGs10wFrb9N4vXpf1fTNrxKPXW
SPo/uGItbHTU0rWc2/EffBfm574USO/oCj8Zo9zoCzoEGueCOItwmSK3N3MmlOUkBnOUgmE+V4Ji
ti6x5+dCElC4Jmafr8jXL7ArCVXK/dZkB+GCXLyjuksk/iwrNwGWBWimYIshXVDU/enNUOlXOD+u
VRkPz3AcafilQOfSbmxn1zMGT85OGYiwbDNsp78NRrwSeK5lQHhT9MMNA0fdrvmVLb7FMoZN4ce8
5cx6swZZm3Ade6Acb5ezADmCWLKleVckHo+oJfaocZZrs77GKrfL4tHlATJRT5lokzwYksw6t2cN
NciE5c7fB0qsirz8BnMqhJSStMyjhGpsuEayY2/M5b1+X1Et5uxVmv5mhslSgt/PBif26HMoGvnK
kyJ+dr0DtcwfcggY/JLkjCy/nSbqUw6zfEV+KMfLOLREPt5067Q14VGMcPlDuIEpkD0sT7gL3hn4
RHCmmiByyIQ98FNpwmMzcUijpun/RWiw+/M+PoEY9ekXfuiATxasAfwOso/Wajv1ca8hDm56D5M5
SX6LDOLUsNabJdReYnfUEspi6avvLtRphwt5r3QIqVSRCp9o1j/vqU206UMxXPbtIBroxhD4nZFO
WFcY1VJO94RMLjuXTmKxAOrZfURVzgj16PbzIYjtuRK9vfpIUl7Gf8LI9T4sVgDNYGMj4atabag1
xogblmCyqMWcl/mTmDe5zyMY3XfnmTMJy3fujEATiNF0D5LVw+qKBc16W7LPxKfMQT4+xBnuQQHY
9U5bCNl9tu6HPHYB3073LGSFpAUl4hMmy9BeYGENfFwNUqUjJgQckEbqy3c6KoQhIK0EzF4IfLNr
ePqMGCKm+66nEDUDS5DSuH49mA/wUWywk1HHj2QKjw8Kd+yiAytYX+sGy0K8+jULF07sQmKk1vdT
CkDeRPjA5tcaP+gihJRnpK2+O2Ch+VGyTx+nh3RxWYqhjiHL1fi60Un+9E2JowY0xd8SiNLXEJ8s
RO7f6xtk0DfLx4sxKGQeBR+aKoePcOC8y1d5+mVoFfA90pcqtWliZ0Q5FNVm5z5rCHFM/XDvKQQx
cCSK9D6HWrkv6xu8vvA4jLmAE6xTKls91jjd6D7o5SxX+DM0IDH9e6sY5ewkHvIREv8IYqDW4dHA
InGkP6NffcRrdCfq0OvpDJ3IqRwiGDMzFSRNUU3tBsDv2nTWJrEFgP/h8OS8z1U6BvHsWYko+ICP
A0UPY78iSlqguO8HNHY4J2mgLcc9aKJP/vxQQtPLa675lpRQ1zOnHaG+KcZWsanZ+huGVQOI0kcc
0gp078Tv4Vwq7kKYyu8/FWPhFhm7kMyq5gqmK/LXJZe8IqJTSigOQJ718oydYjfk6wala7Mn9MUB
/5t/2PupzvF+FMp4gVG2B7vgqN06BCy8m5qLLDoFKKQLAOeTWDrXJKVmliGD1j6DtPYe9Vyu3hIb
HVn/UnPMUXIX6RkW1Jw0SVwjEQAQ16ZuJcS7gqtwlsgM14vZ43Dn1ZZYpuPIazKy5Gh/IfaHE318
fmaIapuvpadWiHkKoPUcq4bcGwHleJOEdNY/3E5DOoyrzpUKZEzsYNofp9ub+T9BfCuX9cQ5oShd
TKy5dTnOgHfpZ5Jb8NNNXpopcMYhxDuS91K+Xwh1xCbJPoBGgzwSTQpYBkf6PHH2ngQQNGlgyjy2
iKWgwrtNd6H1dOQLmmp8D0nKjDeinTPSeyYtLRFUjCXyKpl6BGJoylN/rUuoE36c8Ixe9fr50Nm1
lrRi9eidBIh2ixL5Zmb/wGBUqkbhp2TUUkvD/jF/xSji90UuYDERJt3EoIE20QXkuKkEkyAh09py
bTsh6oBtgDdDpXlFw1QLebOPgg5FjS46Cxo33URAuT4hRzBt54lKsr1YhN3AMKcttwUAmXOLKZmo
2NHBDHSda97VyNuGfQjXCq+gXHI1cctx4WfsGk/xlog27DBW3USufcqu1Nv/WRrU4Y5rXm3A6kR/
Dv9u7kaj0zJXf0quJO+xKH1iQjstClVtgazwfHEH/fTx/ECTSJD80NgJyZeTSOFyIJrGPdHouQB3
Am+JBhKeccQqkE7PnQLV40UxClJ3J9Ty/ENcwqroVgyr2ZVktPIolQXVoSOVe45+W6ijYbzSDCHe
wa3oMK1i0jt9GEn5zHQBUWmytTS9m2w7NQNwK/DbbLy/SWIN9pkH6dmMlsYRwvGRtndvytUXDtZY
rrLbKsA6laaXC8aD2VowBn1i5XobxDALSKbDckAJpOVoIaIOglUiDCQeuYgr+kfnRiDcc0I/I5eG
3f+yO/c38FWTlnX4J2Y7QPsckGWtrAWpNIPGHDoiSGlPDarFmwUcUswthcPrr8DcoGnJOLgl11gX
iK4obvcMa8A4/deBd89hjZ0hJQj/mu0DVFuwfP24CNgv9VdLXBVmWP5w2w4m/9CkkJ29CLyMSZGk
nxGQlOnuD5IF8Fe44FStd89rJDPYQhab11mfkkp6IqKv+u00r9M8vm2dtO4PD+swWRWA8/uD8iKu
CdJPD2LG13Kbfy0RtU0b/Y9W4WVJERXd8eAhwdwYlahHTubeIJZAp529440MRw9qGHRYlKBsjQWO
33r7nhcwWq+CxEK6raeod49AHimTe6PzDPVfosCt/cNnt7eRquBHTBZLpnDduWbPrjh1e/Yu9YBp
IVftlcvJmROzRCMK3QwNU/cNhGO9U/9uuacmONTEh/5lK+XxIVpl0wcdolyBnz5T5fENGWPlpRno
qKMLyBQEqPkIUTAayRpWMO4X3V4TtQfMA1WLO8BMEfKgu57QdgwAaSQkPweaALrGEee2+B+7K+m0
BahV1kQwB4syXh9T0OGC8BuKcFPnlo4rZLCu5JBgOp+EhJLeX5x6o40/nvUXnDmoWFaiY1roL3Sh
87JpT+sc7yfghU31Hjxe17QSxE+fpc5y7t3h13LXl8SnWYj2lDiDIe5dR5sh67WtWbu+li0LRwU+
KyHackp7BZsBq/o/eXL4lQlfwWLLDR3Rp6rxYbjQrtnKE5H+zZWYH+scGHaDKelHqpaPBnG3WbC4
LJ5z3xWpAT7w3GHGQKlSWKDONXfoIU/rgx1B6T08AewtKMLS54iK0i0khub6lu5IgWy8OodvoElt
sKqsR9HxpXHm953rF3bbfl8z7UkKfI6P6ba4bYCbOPpvcF9dbRv5arzU2nS3RkhDdZL/djX4XEtD
3UnWIh3RHrsG+m6szBsn9ZljShoDvEiftaFhW5iI8rYgATUZYXSAVKb9/nDAto7z9kjDYgCLEau8
h9Ob9k29vjw7ShCVMrQw6Am9y99B3ZpV/sBIeOS1mwh3duZ8KCSaOSEBIDXL1P6hjYDMG0AxbI0M
zJeh4nv4yiuQpESdqCzFuSAplFIqO3RqxXAfIxIWBsn0T6K/VLm98QGgAOXTlDT+RNx3F/YuVwZr
zp7S6ZwjeRdr3GrabFce6u4cksHCpjKRr+6h4nogbGy9adnwUakKQHdSW+gjvX0/prf7lGvmQidU
ekTZPhByJ6oENoHZlpgr8dcRe1bCMHbBhYflLwHO75tNGMEjMsBlZfj1o23/zR2kgfs8eI8KQ3Ag
vwndBDq62dvd+LTr3rrGcpnFDqdMz3ALtg6NMY4otx+Jn2Jvlo3p/hzPyRPKkCCNeBqWEhNr8uFw
0z5DFL5Mbqi1n2wSf8zmLvAdvSd1WsahqJOEbE2bWPlj+jMjaVLzKZZodgQvKfwi8tblOAjmqUih
pLOhDEd/NajMuz82Dw3szb0z3znkErs/0ZvBvgQRJZCEV597ggyZ+wz+o7iNdLJXlFFjB0QUGeKp
+9tfjU4E+9Sf4m+S8IzJ57xqE1DpwN9Bcqu+OLwHV6QK8Yp2ICfbVmrvCtUpJAy9CPsd25tKI9VZ
IT1ZNY4YgiDdMkJ/wajfTKlo8G77d5N5KkRBACkvj9ztqUg/OTj8sO3tUVBm6tDr8L4mbltuf6yU
/cDm7cIG5wmRMSK6+XHIoJ3F7DJxy+gg3zxJE73ScYml/Jq0DxF08e1uNVgTvfYMj/tQ5nRsbE7T
VGY59wDUNJXpg3NiOvF1YOx3Wm3h7ir+CfqRWM/Ug3ed2MIc/jyJlSwIJk67GjO/HgU67bOhosXB
RjSfNwRK7ydMDMergMGiMQBQnFK1vgDH0bwEne/AV8heqUJZmbRGCKPQaAWOKQ2K/lFXKUbPXqVZ
olEb25K6R+qLJUV6GhtByyR399mr3g2AnfydlRbLd3aZyhlk2C0z2BvPnslqdxww3tYvj0mwzI7j
Czl9al2S8ntTrTGj1skJ3GuaRGb7OpK/26C2KOD2oW1Hg/s5CJtcFJQ1oi/yblCOO8agHd2GZIh1
2QDPOJxnEKQuPlhQRxnbaTU9YeD1gC3B2VgdxcO0j95KEhmXSVheSZPEFO0Ain8P3WWpoz4E+b/e
VO+lf+Teomde/YqQyfHc3sQfjCdAGNKvRRqu9c3tnewZ1K/Gkmwus6gmEeRz886wtNm3y4CV65jH
CdQ694VG6jEJY7Ht3/9i3z2GLMBJOYeu6XJKXcfFbBhTyxzvYcsK6zSngeeoNQvGsE2eJwcfex5g
6t4fwcgyHbB3o1euwPah09pvK7vR8/k2HxU5K9o3S3p+DK2eytKTLWT6J6QypnT4jPfaSUo8vvgr
cpu7iwe56kFemUYfWdGvHlgJa7WppfWo4G84NsQr3U4iYWZdcmLqVPrXPAiL/Ij6ZEgjHEGY0v/n
yK7TG6OVCaLNuGOMNisVqI0hi5H7jwzFuxMUXlyKBH72DIvuA45JBFB+8MdsfPQzfNEij9M0oPK/
NnZiP1L4Na/ny2jOYMD3+YwDjIm9eQ99Lz8+0Q0k2Dfx5NCsBrQtuDcd7FYC0oZn5uJr06OHs/Mp
yzHV3dOhoOecE5UAwyHPpmvJ8KzCwDFQtgZJLTY6ROHadz59CXsPkmUT+X15ijaOoroH8T9D2s/f
t51dlhOv6eh+zgRVSNucFxl+Lzg/svzEupdcLqMcqrHzkHy60ozsHkquBZiW2GDHFxQm+VHBVXm1
BCcSv9qTnTGONVmMdFgm03rERS4iMfkYYnwgpc09Rr4CZR6apVGzIoujc6Bnd8bZHsKKqTkKy8H/
cLb7DgnwyJ80RfpZMErBxI2MAfZJxap5cBqgaKJwj658DuuA5CnL511DN6Vthlhws2wRsxw97TA9
PIHLzi76wYZlPejCaOOMhmUh5wX37zOK9U2q0cYP6CpZmAHCCcKKYTq4FDqoePYzF3KPOrf/IOUC
Mo4+6SC78NKH6dxmSI3TkZjKAC39a1ep/dVyS0HJeMvPZne+5zj6pGX41dl0b4l/AFoFzXl6KAlJ
H3uU+SOMZTgSeG496rk/OOEomEq5KuSweUTv2kg68oEcx/i/ZKZtob6fikiJZh+wTu6henifipkz
13FtSwN8tx7vb6sa/xk36ItZrGvBijyBIEZwmVwVwC4ha8Oo9OmUnO0AKpSpGuAaQ0YbNYDYbRZ3
+k/qYOtwcUOYI7q7r+/X0P4ysuQ2/Mjj661ZCp31YFFC2J3RRcRF62DXCTcKe017xfawVAZtjvpV
vkb88HLaaAwjjDKgeQvkEPogCJUXyUGiyhy8PJuYzIEfd+z/24ncU89/U7k35XXeuUXbvxxVo51T
gkMK7narSaTT9KSVV21TZRW316K4lerANXS8Oayncrfk6mEnWfXEFDUklqfuW0ie93IZAgme0Btw
IBGOKPxV83BkHNpg8aYjFw7K7wteDQYZF3yF+oJwuqotecBPKjkmRXIrvWY9HcH3G0fowZkMd27y
NFRRqnR0q/PMbYpdO3FJoWi4Kd7InGAurCj5GFS10hl8dJC/Gm1dRijioN1xtZvznoQokUXLdJJC
50DJY62ZoMcL3E/HahBZqMQLZk3EcR7YwiVyU9xo5Wz+BwTBftUIwVPHPgsK+dYlzXanXWKKvBaS
QWAkxi4GJ0WPnWFANzToqjKf0nc5s6S9jUFfKZ9pJ0kzg/Hd6EHaCT8uJq6FveGjAaPecBpk7mxN
4UUUf7DQeWAtN99R9hrsDrCp4lA10DkxYpZgetYQVeg9NVMQJGMkKebFGxRfik573fxP57vDxjZ7
QgcC8aK4x2z0Q7avU8FZ1Ufhm9XeRVj4JRLxzmVx45aB86KwsH+yL/vJXQYFr6oWX4lxCue5qKMJ
vgIfEpEUUxQ6P6fWrVANs3iJNPsUOmEIOLR3vfTBKWadD1fq43x0fMKHBhOv+T1rHR6JUKFI053V
b6fbRe4wZQe+gcI/MQbTdwBp42OPcEMkTShufNavur5/xIYYBVQUwFVdet7CRqjHP6qNGBrQuS/o
/eDThv4sMwCPjmsbKkTUX1nnosYVCryHJia4gKHljC9AD1KEUKScWQq6tlYyY9apLQmmRtmXdV+s
7Qu71pI03mHus39HK/nSM06rVc0oTruu67wm9+hL5t5TRyz4C1dWpH5/LPoG4bhHnCqMghztsH6X
BA93uvKV6+vRS6SwU2gPxJ6GKprj1oSJhDobKFZQhCY9PqP/Era+Dd+EXQCWjszfbwD9ykOxxJcA
J8btb5EmEGC0nEvDpMJqs3uIkmSs4axt6NA5vP+gMGOUbZnmKDp2M7zLILHgCnu0GCZD1IOa5Wre
I+9wWopp2fze6CHjZc/r3Pjne0FkwF+FzxdoPe3XTxEtXyaGbfdGLrwh6xKyLnzh6d8XhELFdn0t
Aj2mklkzZl7dynkt721ihW1uZI2LU0hFB+wvAveKA22c4Pt2wvGP604V29kOOZkM63yGSMqYmLD1
mww2InxSrE0707JR8uvBEAXZZ6M5hmIpbujevfERMAVa4hZF+UW26u2JbOvE6A7AzbWlO6uCDs6L
RjF+Y+OmhgFncfC3paEEjKcRtbBLdz9okhTUVYvcJMHZuwECgYZLqmE+E1H1jcMzsvvXSeawroxV
jPb2Trl9+PT7+XIZs4CFglDsBP0H6NvAoZU6p3PHe86yWKMTsm7ivK/XGFqDOX4c394fNr0iQRXX
zyIFX7twLuIS0d4msks+jYWUeAv84jbfojeRo08bO4E9t02FAi1F/z+q9vtpI7A7BxTKndYa1UyA
15cePe1werrHRqT14+272e5fJTK0Tpxg5rjJ8Hqnurl9oqnfHaqjD7dFOU6tmt7tRcSDOANA1uKZ
u/jNjAHceMA1q29G362pxJLrB03ZmbFMqnRLaw/o+MllBKAzknEB4jF+JFO1cRvehaQxqA1ywkgS
ddaCSBIrjAkhsPYycsePvhTAAB/3sVwlCRZS6QN/czh3L0HzEax0hz51uiDi1HGElOaArIMzF8QK
DvE8Ib+Ky0vouHAm06RECpUj69UDkW774Q0TzLaivzYnuBQGuq2GkEDfSYHBLR4x2WS/VaPqSuc4
jkUDVr444DGhYQZXcCXDg8kGsoYJKbgF+wPmwQVnp8kWEPuy+wfkdawGx4y38EV11qoE0DTEJuJ1
9lz9hJwa+guWtj/TWxruA4xez0VusG5R/IrPurO10TTn4Xww45QY3+QysKlWM9zv33jjLB4zA5NU
rIr3spPoJQL+F8BtAw7Pf8u/MY6++cSPd3AMQPBDDkgKiCGGbDIyNKR1KFOO/Tsw8gfQlpI7WwHN
UlCNGu/ItoEQE+IsVnnjRobVJiC/yP6FYaoW21JXg4shovq3Cm9QFL0buWRr+JvIi2SGX0XqRj8h
PFg0BNjjs/KEO9RIyfO31SAu5m34duJ/P75ZjmBK/1sBUWKQ13DMIS2rrf3GP70g/+AukFIy24sB
QT0tti19BCUE46ytEpD5TYXlm0unVm5HQrz5Wq4uxUIEaWYf/tvvcvoXYbsUvbmZ5pdA5Ti9nkZm
S1BncMJUig3wSA333rORYIVDH2I9FFp2aQJFioCNYr5Zyq6CHExRc4ZF9kIHisv02Fw2X/Wqmjhn
vLeqENZ9noAytiOCMbhzih+tXGfvM1ghfejQVM84xl9vpmZKOUZR4KU5VwB5UxotZ11Geq+8MQSh
TqKrMvYrxbutWec21GRVU5vv1XSXr4lvWntTi09kJ2RjD3saoGETFXBsvhkl8UPj4BXfL/EgTLMx
XN6EMaRUkpcmCI+efqN0UxhjQ5YqBeWIyRr+RTtG0mcNYtx2wyRyiBA7SudpTl9HRQlEeazYUa54
43ynGEcDiRXa+K3F026LtqzeHC9awQnVvf7LFifvwe7eTh/4jG/dUqHncE9WkX+Mj9t2c6flUcnW
98iId1fRBSnqxWLxp1et0OM41js8l7uhmsqEbkWQbs0Su+W0JgRIPaAku9HxlmLldVr1JJxq5vfr
IMAUWU5BsIWkD4NmX10r7JT45HnqGhVdXwR20dI+8zJW+lBByv/hR6guYpeI5ClX+Pzc0z2WEqX2
IqNeyKxaYjYBXvCnSy17YiTO//lWon6htLpEAEry/bS9XoTvjF3aTGhJtn1dNiKe9Q2wwA6+ggNA
2Z/2qZdCkbJz+/rgBDq7GirBqUhXfHhqjAhz18ChL9Dx97ZW4QheepnH06Soms5ySYkwv/SpF9GE
OrIef26m2fCj/zKmLj6dJqfqsKD8/z6GuhqSO2ZW8bm23nwf+zLIyZn+Tjom7RwH8pFQvmiwPU3P
N3tjtTBCa2YndwdV9xD7Rb09fqZDnsLh87bR7Q8+IABDHtiXaBFwegcZbET38mala0kZNL2KO4h7
Ym1+KYZ3vUWRIRXaRDDS7nyl5l9QUgGDOQzpqj7yYCA6ayyu42a28hSmMq43uAHBeWH5+8Kp0q8O
ajqZ/9ZXh4JCi48sqaB/PMU4JA/DMQENjkzDYo34MgIdmLtS3hsTLA6jhqVCb1WGGK99XUTLkryF
VCQKi+nb9cpQzlyr+LJpBVm/15uhBiZ0kEMNhAVZzbz6YUeWK0p38ycgumY6nCTFLz2uGWzYkDpZ
fxiSbJ5azAEFhEwJc3QOaRRbeP3PV7yL80jUzfFjhQjty9DCDd7uEgJykmPt0Cpw+x6zen2w0Jwi
ZV8ImT+QdFiaVtStDt0CYwNIjCrjl20aDHajTA1XttTj3TIxYPTEV+Hpv9F8/3cVWMn1+mTHVUZa
8zQoW94BJQmzR0+8cu5AF6dxCuNN18EkKta6lQCcHCITAft+3q+09kZGc36ABLJcZ0eVUg9noJ1a
YuWfHSvwo07cIpqNlp/PXALPshIgpAZpoOr3gROnpBQe8JIZ7RU14B2LOkD31E7I8sjKhLgEGPLM
hzZM+U3xgQj1zEDMxUMYFRs1iThpmSvs1O3rzJ5RA8AaSB9eX5FbaNf+MPBHwC5XOXlVDBfuVZ7S
NPcq9F7tL8YMqIBSFvOsw25KXLoqjG6QlKCdGm01PKclB/W5bhVqY7nffaXmMfNo20QTDBh0aDZn
K1eeqjq7mes6yTUzsOVX2o9O6dH1fuWqkDbVLbKlp1qh1cjQ8mU3+oWPA9NT9WCEL7q5pzJSVQOH
i/ZdTCO5UuPM6FzzHV5E0nUUYBwEIVNgcIkvyK8uoax7KaG6AjSAqjm8I5E84wBZqAS3VLFMlr0t
JhbwfifAQON5LRxw5Ozz26HREynzoSFuzwebcpxzot9PPLx8Mmpxbtk540U9kTdtYts2Js4saf62
nLaBv4H/yyGW/28nhsjGnLgpH72/+vTMm6a+RGocytiSvBv1tlPriMDc3E7YbNF8qJf4m+3CvdsF
nmLxX9vdfOQBkLRIPbvWsXq2fibdKv9Uu5ZFAtsdsOsFnCrL3ixu+h2rmEvxQx74qTl7ehpFY6R6
xcbAPJDSHcd2E0G7ESNu9w3F7sc2A9WSNZkFwC35jNWf+lUd4N3xVfF2aSuXBrk4tsgjVpxG6LF+
+eW+vb4uzHDd7wNr6jCQ1MNXqzKqr9Y9Ywt1hIXSUVVCfAmWSln7/LRo/ZIB6ZpbBRzqU7SCK2aX
XmnOqCPZ9tLdmH+ds9j8Fj8r+KZD0dg1QvagGyXxVATVfEOgKHByxvuRYqAyl15wgcKSf+wpjNz5
Mj9zU7xFOHWNwsj65JWMkWuNJSK74wnGi+bkM3PMUJKT6/OoViUctNy+cwVsjxUCgpysaHjkPHfS
XRKgYLKSIVJ9NqK6KvGqiZI7T1MS5JsmnnKhdy2I8Bajb3JF28YCcFKfk3JurZwaM0XpK58O6fkU
Km1AGJCwxoxsvzLubgM33xRf262RuEHfGyUh5eYGiqk7kXsxNmbGzWwjW78YO13PLDsR0veEUwoc
nDk4j8rbDSWuY1digiC7siATmXukajhR6zoaW3jDIyQrR8D+hsLqOViA9dxEIimMemxupZk1Fc3a
yQLCsjfmUjkITink//kw8eSHHjgl/X4aLr+CkObwlnYi2J2Q7pxyUClFZIOYqKIqPiIj4YFJlJUO
PhNew+q2TIp/KYoLTu7UkIfG7pXwHQFl9/Re/gZjZ5M4iRKasNakao58/IHkSBnRzxgFlCGlvbuC
uD0pB1pKQkoeqPX4zxLUhX4Zyz6JrzX+sX2/PtecmBegTQx4JznRa6RM2PUoCzIq0vV4GNxTn9H+
Go33gIMEQSkVvl6qY7q9O972cJUAkNJJNCxUpa8D8qJhEhenMHhYxuv1FMRLIEAV+k6qaKk9KhBm
vVpOjF9276jSd9wp979DS3eYoJA7+3xUAeP154CjLnT5NH+yzi8dc5WjLbAn+eF56oKJ+jKlgHMP
KUf3YM7j+vFKBjXJYukf1yauo6vKyeRI6tx1Adz1Pp1uPkwB1AjvbC3zaehwqwwce/evQBAaZM0a
XO9q/q9er57eteytwBwjLlTqBjzAv8Erj45JMi4U/O/KeelT6cllyIz6HfZ49yKOWIVjGEtz9Izv
loLgVUiaMi9cphqW+Y5CpRC3kOczhQ5UClQuYTFCpOPSbEH18N8r5vY2iWSg/1h9/g3f5qRJk2SJ
pC2nLFEibiZRne5RTO77Fco5otf83p4xrnfobEEYZZQFpCtxxSDAGGv4+8O8cEfsNKcgfSwA3eD8
SZoKng8HCXeRK6F361z6OlDX1yTk5l06CsyuFXQ8mx3T0jNRMPGg8uaqJMgrFv0zx4ZbDIkQqKDr
oNyZJW1J3mdkl1l0htFtL+iLJlr9GM/dialHZcXNb2OIl2RmBulC5hcpxDykwgUWBdo/0Z9ATAwN
LN/l5/QHsVBg4BBbrzNlM/+AFof/76B8StDx58shwyRFq17+h4lfFqpUqzSAeWGx9av8V0uXhrMU
nAqMXA3znXJNhRRhyBpzdMxTe1Ds3av72TTVmjJTDGYHbB1ZjWpwyzP78WZvAfUL1xH5PATJxj+A
eE9wrcroTy6EPFLAN6y6VdrcqQOzRtduBL24AY1ii90rU06aipNhjzUr+4WrOqiYgoCXVYgFl/+S
ID10DCEmfw7Q5dzP6r7nBneXHE3x/ca/D+Dy9ARcWN/oMe/VlfCQ9ugaACz9oW1SMYyOKC9+yKuo
/8JIDU4Jrv/Iml/m8hZHOO/3Mso9tgC15EQPQ/sO/Ww2FffWFr5+EmCyHpiqEhsJR9i15U4aQK7v
QxjjR7vf89VRqRT4HU3b9C30shtZR2h5HEmLRsMhcEoBf1J537eguIp1indXjyfQwd+Aa0cFPAsY
YRuYRyHHdreruo7OsX0RSQylC0AXFvhMjw22UPppNaw0rIXfBK25eUbPdbu7AaGS/dSBj1jGLRkw
2aKZ8lIU2XWKgOT909rB4LPzNvaayNxOeQXTWq+sgBII8wu+YVZ3avFnfcXpyBU4TghiBU1vhs6Q
/cbErLlS7Rdqe7PF4qFyusMZNhKlxRIP/AhTJwQI4DTsIlJuQORfEZLvc66W1tsil/gCN4q63KLO
yUrdrLre+zLfMdn/HhjcqKKIaxjigQ52766RwSxnXunoMpG4IS0VtxHkV8tSjQb2jQS13w+a4Nbb
8FY8aA+wGuRv1a4WhHCJGhCP3ZBC+Iuo0ISenPlDn3ieEAqvSkDaKJeiUG3PES9BzBOjK+gK7uqx
Pe9l6U/+RhUM5svcP2gWYV5YFTdumF7wC/fj8vNkp7MR9yAb1f9i5ZX7B3U2dhIx3UKpe8GIgMIx
DFs4ALZTOWhAxHXkAHXM21iSn94OXrZFB6FVFK5A96cpHOoYbH2pORav1l3W9hJJiTrUb9gSbpFI
jfD1o4oX/0QljRaBAlKH8sXMwl+ceaUQpnX7fqZqziSaWy6u5lgD7w9skGycKTQVl654ATgOSFcN
cxb3ILvXGpElyMtkhU3TFPSraZ6ExwYMdkRMEMDGkRuWj2SJCzER9IqrHBp87VdA4bxvNmmpFwPd
1OPP8gld6C02wNNS4pi4nsZWTjKPrhZ9h13l8uhQJH4x5UXZAnR+l1A1+DsadTGOLGjFaneEaobL
54GiYqzaJlmjj1i2aE4IoX7E+g8kMyd0Psqi+yaN4ob/Fk7tWFr3fu4XBor2qBxTQ1xV9UFTiKzA
G856aOF9S+zOxLVJ8teZ52Bd4cMU0AqamaRQEgrotqup1Oqir8Yg8GSjVorQyo2M8pgFmtolCdAi
D8ZQnF9QJnAOqq/A4Xzja1pNgsrRz0IQSOezDE66HAsIvYbWsGLf4GnV+DDAZGBGg5+gZqL6LXzQ
vCZPHil7i8+FuUPHMYDFrSeKuRtvxNQ9UplhddpjvJjOwz4wGeqGwExHcFrr0KWPhRMKgLd2L9ys
8ThzvSrOnFUbkbnMaYoEoMEqdbtLK5pjZhctKLsRLaOqZIeZL0dWEegGxxcotR8+6LopVPY0qfI8
6ZSG1LpJ3buDyjN/uxFld5zTa9KXdYNz9NNQR9RnW8nB4ap7cZAYhUIeN+/sMwlzZS9R9hBVYsOd
cfVz164YnU0jg0zhU09nGefvqX0WF5HakQtvy1VSHPeZrP483661Os67XTkPd/e23AnJikOAWAey
eQ6u1dm1v4dmpgQYq/QzIzGnGlpX4ReuN3c+5xTmwhRnmHHXzYkF6JyRzyJIjUalVBCaYDRqaZ1z
ML8huRSb9VPFjIxGNBy6liYNWGkJtBZPSC865zQUvd+ZG6jbCuO03IiMHf14m7XqVS2JVzLdPR4X
mELPWA/DjVjC0eEIyyxRg8pFtJ4hxv/bWeaMjbtulvEWC2a5t6kcQYotDfG/liZW0/SzoGv16Prz
0jzdBKK99RRGbpzemIOxaCGn9mWOsBPlfHBPKcnsMbKvnAACHl/vqho0aB9nu9LpZzCwWj6LI8BD
n7GvnXJiKUz2aFR1DmqQRAPed4foZyM855ExpzgcVIBC4umqrjvHqvhYTk0XoSDMPrDGKmXfoCh7
P3X8PRRuX7CdlZxvd7HNsyOhROeoDVCdnnnyvzbxV533Tjc4roRn9FfgQ03xWlfHIebzPCiYTbcZ
+xR0UOenj72w0UFm4Sf5XRP0VhL2//E7R+uDsmZ6GBxdFUwnSOE6BSwDMvL/R6PSzSxpAalTerOX
FzBtOBKbFmVn3KCc8fB//U5lMIwgvcjTTqWkuPbcJ9/KVXqO1RWpUrO6ckEorGyIL9IfrK3dzDgh
IZx/h0C+1uTgvFzlcrFOJ2jc+/fzPnjueJI7EzfzNrP1pzspZWTODKk/DI+TSJ1jqPDkN8fmVwih
HLmGD3wDV6gRo7JdqcgPyfYZ+DAyNMdNnYyIU6rIOp2apbks89mPkwiTWATECv3h0kwblnr5yA06
EyrIp0DmBCkQrMP6NyxbdozywviH0xVlDoH3cY/s4h/NjDspbQdc9Jrvibb2/O9ceEV1M3NlV2vX
krWghy4CFz9P4Rhruz6e5jQzfUTgaCvYElZkXdK1fpdFWr8w7LCxydv0T8NTu0fIuniqEQZhDN9w
upsnPbGAaruKteZrJzbS/ZnFqWu+ihCK0cU+GfIIe9T8Ygfl+o0K1Hh4xJUDxtYFSrjA7mHTWZ+5
XzF6q86728knNPBi2pxvkJsddEcWWRlO1OjtuVwQOTE0uoMGJRSZENmGvUwNmw7pOfQnFw525E0B
lA/1agWYMsQEVWOWaXUpJADQvDAPIPFwNYSlYRhvVGz3Nc42EIJ12mVFRnJPA05ntWlewa78b3nU
t/bXCZzC+QIVJOyu84gyElDa1gmMZ6jPWQjj6jBe03HV2spPLMXLX5qtw++A1JqmeBNhapoMLZ7v
nbd2z7zKARgvT073zQaQOleUdlxmGLd7nc5glYoGwLKuNrs9VO1D2cF5CJre+ljs6ir+wwk75v0P
zugph8HTHZnnelDpnpLIIzjfoJVi4GjEm54QMcerOMCSYGf+0SogqASYj967e5+Iukhve+vEpn+V
AaSOzMgDM14Ly6WGA7bwQ+LrQa/rd43IorfJNrJt2bc1Bs5Gq+AmkVH34i1Ow58NHH0eOIOft+2b
1+OtgAC97YQyiDDYerMG4zO6TzJ+Ei+CC36gS9LN62/YhDtChpjQY7fRGj+CR87nwhqPNHrspHnt
ZJr90J8zeJZhJWBGsKnzk0bM/ZCxOql4oF7Q7AYz6rxXVqSTFDQum88YdDOKCocvrbx1Py7tC9OI
nwAcObZBaRE8ztXU+kPrHXeYIJ3Ga9C0iGCB8eQTxRzod6n1tsZY2Icp3Gymku3k441SeDQeoNWL
hzqek2nofarZj40MF6lUbVIx/VtushKFrpnpsmIyt6HfQzmPZ96irQcXopbaDMfaJuYziZxSTeql
628A9JuxUyYByrtFN4yJVEyx+DOoktZ373nkVP4gvsRC0b7x94gj03tqbSeZq6WIEFrp598jWDoU
Ic0/HO1JOXIytjLbyzhdpsG68qUgHhVHjd1svX/6Mnv7BMW1aWZdk4yFUB4YFpvkMHoWq91BD3qm
qzCM4lzW5fWJGnB1GapstSlqTEbjmbHA2NTVv1gP9LiXvnGlwDJfnK+D2th9O3c2iIiOor7ZO+1r
lblTCuCIfiBTl6tUwLeydFhl+uICvXR1u6a75bJTq45irCE8OSa3fpPnCFVGMTFaSw+w3UGkiUCV
rjqo2TWYXNZHVpoXLNtFPOQ5FYvOEj6YFZLWcbvF+MNnT1uFcNdQRdFuNtucFAjaccqp3Oskb+su
MJEcKr5LvxidWR3gZGEDYUj7iHm1CXTOYEYdNu4KQfuNHFL3XbrIc5dR/ZyrVna1cWuhgplD7x2I
nKny4FKFHWcircvwlFpmFsrmzNWXngQxPqJiyD/+2WhKXKTPMuzf7xQtHKlO25k+VAbLnRuBmfhF
FH2SQEKrda2oyJwvklE/VYbB5HxexXs0avBLzoKLrje0WQm7RwzdBcYdXbRvu526IMeuYLhVkq74
gNaV3GwN6AwLTKDl3EXMDJ1j7A10NGs94qP1qMBgdtQm+gyk++/LxyGfrcTEcE4/jessyFM8+xDg
H4gyvQJ1Ee+582CAT5fReC1F4wEsSfbtwmDUEQa+JXxaancdxN9jAKtVQMZrREPphI21AtvqaRks
/9XPXHPcfRZVJIyddYdIh4u2EqQVTk4WA7n82faLW/TvhFPysJU37hRE+YMGxZUyz/wAv5n65Pwm
yc/JtGkvUqUQEwsoe1zUgyXESN0c7YmRm6uHoMWBHX9EXwQh/IBCDYNl9FYi28sQIaEP17/VBDUR
xLSiujfRva9qdiS7KUZeagzjlr7uYJor3p5OMiVQrFg/hsa4R/pp6OY1GHofQRL27LQ4J5Ex2INq
PV2KAhd5SWh6U5y1c9aE/OKK8dNFEdxVWTUvgI1K/3K8uf0eb80SpvMpGZzJxLKqNG8ws3QluhF8
oerr20WaMhyuq+ezChXSvxvcv5KWNaXXGcqC7H70rmpzf0F68FxY2yWCxNUpIA0B0vQy3OTq4vs+
Fsr3lXbxIsc1T7+bK1JIz/ZtyglX6WKk9b7/p86NuYAt/5eSWLjgIkvgG/8MOa1TRbyyO6oHKmev
AXgVbKFLnyPmC+O1WVgwEtAMG0yZd2k8i3BaerjyrHfeWaOgZWHEA1illMgGHUAHBqo3gk6BM2qJ
zXw2EHbCLnVosdmlkMGW6uu3eAH32xJE79sWsZt81lQgUBQaZ5B4rmfzoDQ9jgRY0Z3iOJzJPIKS
5yhBQUPN0dab0CylCLekg+vARWLQUxNTjesulbVlJucRWSrE1JNtpDkU2y9kedFkgtTcRBT1ebP5
NdayQrcTk78pzoZ0RB7vvhmwTlwDbgtfS6oegD6syIlc4524nFCDmsTsRGk55k7w8y2JGfPu//6a
j/rND8lGT6hoslC2EehjwwJ3saw5kYjTilptj0zlJTRVOAV4Tx87rwxqVZv3K1D37I7vQQ83tqB2
yhKGHBIEe+AqosoAnKTn63r5oEZ69J9uHDb1gXuzmjl8DRkOalow2TkFARtZt0G+6CO9MLJRJBSD
X6zDE28tAaxfj+XSpTynrw7hN5Brcv+sLBg7AD020JpOOMcSPcEhcchkZ0wEh2Xv1eSIdKaCZXWx
jn5iV9Fr6i1xtcQREaSgFiNdMdVDJu3xrzY+t5RZpm6mWCMBSUXzb2vyrnkvnYshzpM68r2dh1bU
n34lSy2J7UfyaqBR66wcTSAgV3fbUx9+7ixWtW2ZLxbzrx63hdx1RXB7bYItRzUOgb4PhScvOPcY
fyiCrUzH86yWSaFuyWf3CRAPU17PGE+jNzwrLuiGqTXB7epSX4x5z67thyoAfNpG/JwQ3gPHk1Fa
vKOH9KeBHHznTvIRqlpmIP5yuO37GVuNuhLAK3Xr7AwOwIn1qodooJ+xDbPtqVUH2aMy5S4NuXQ4
wsRd6TeaNOh+ZVUlhx/tVio5URLNBCt4L0+kzMIAx25k6T7oy7ABqFhO4BimgQLkuuJiSv1TqaY9
/QzDpzG6rsevbGXWQzKwEhac+XxIMGqvMHASFsa3x0nQhHudMDEhruogU0O03Og4anxF/c+G787t
oekBiMOk9HgrmWUlDuwgm461VqqfiDxtzNWVkhH2YGW/Vr6flxr0serwnY5lMuPBI/v+5sfuMaBO
uX3GZobE6O7I8RhLlR4u47ZHWwMxHn/Rgg7OhLpvHZvxhoKO2k8fGkxTmxWGSJwyja3erBN+OZsi
1i8japimEFAIHhVFJkBJIsHCRv31qWOpF0lj2aJJkRFAmDMwzXVBaMnYFa/UHHYyjptI297pxGPb
N8HREWhRuCqUbI2XYFFp4L0LzR0idW39HJMraqCVedPtiMni4nWtoluzYxxNJF1MXIIkMqHasdGS
kK6EELR0ubUokBsWkJEaWne2jaVeOhxFMSXFCJf9WWEsmleETpX4XkshqwTSwtaoi8PVNZ8Ouzn7
zX0rE3q8cO50cxBvv2AINhDdU/A4D+0tksNaVUJfMmfOvnVp5ntCSVdLYVrtK5vesEopQm6oqULv
M00AiVC18Fpj0/H10fB5/dTIeJw7QrfizwxQtsuTCLXAYVz75MU8JbZZ9ZKLGho+NTTioJBbfqfz
jgaMndnFWxsSbH7xSBwyI7ytjRhlhScnJHlUWm27mnjYNcDHlztFL1S1osNrpT/LhLbPRrtdQyb2
N00eseZ2WcChgjHQJblZLU7Zh5FiU6k/sL41NCLLl2R4NVecGxwF5l4wDwdFlMBiCszRueOjaG1K
fdjYFn0bSX56C1kuDXGpdUwB9+HqaUKVqIh1wHw+L3S2+i3L+WWQIjZGnG2gG9IxBPQU9Swgav6n
j2OuKDZkbxhEMXHPMyC4Mp+ombroy1qz/FxIe9dxZYqNhL1qcDdy9KsGIcDYYIlHFETAs2GQhI/6
qXL6y+bCDhriJ0k+i5DPAlbNqwMeToKd2Q/e6BjbY5Xhk3sMv732VSJ4JnHrzmVYvPgtzTfJj1lc
1L7A2Y6tZuRQaIhpFFvM89SIRQ4YEvGwL8oGZnkVLBM3dn9BWJJOnKs9pRQq/3ECGNEBsdkAsI0r
VxsmUcxmzsUuCfLVqPeDhtgdnVRcp+7uO1Z5QMbhf9Bi2RCWwzlGouscRzlLnZQYpT4ERcxxE1jZ
d5ZSXT3OXoFqv/nb8gkTP1tjmYWTpWks8WoG76vKypq9YVFvnu0MyIY7MVq4OJ3HmLHpJDDI0YK3
Dsj8sEwH67YBhC1rtGvmLIjcHrSgd6PumsyqAkcq0MZvi6UUS3k3GGDtRBZw6tT2f8w2wZAouJ5q
dqmgICPGaFdfR3TYUwLsy+GpGJfzxgKBA8+vEiCr5ABRgcvoBHpXmobYMUeIkztVj6neLXOlcLmS
NXA4iYB/cu+TwDmW2x3V1cMCGCj42beyIqW1G+fSsPQ1PCMusKlmf7+DurdyxC9A+9M16LpGgCfP
VPqA25GfgQd+HfBw+e1XE63wh9vVwrmxCpVqglS7NrFQF76TBuK3etNXfkmQ10Gz+nJgTNZFX1Fc
5c8LzNS14Tt7mTS99HMIH28fLinNz9O6tT7NUuo4+kxIp7d3swMfLnQK9ppK7DAd+c73Zyr4htqQ
a3DSSFRpfMZ9dv4WXY5hzsT3k1d3V1K0Ek1iP42yZYI/eCIs1oBpEYZ9zsjxfDc+Lapa2/xkmw0Q
aRr6y6Cc2qH54cQ9AsTjbFMxEMYFOjhT8PBwv8XOcJqmKmpsE7R+CAYsGfjZjPZoh8OmqqNyy3Ki
f+7xZ5Ao818cbQeu/JqKUYKVN0cy7oLtG9NxGCV8pVSjcvD7JabRwqVRQ/VtWW+Su6g5BHZyjrC1
KGWKlifCpvgZ05NrA7PZ1LT43CGErVksjjOzmBenmbx2FL4aVovx9qiqd3nDi7GtuiYa7kFePu9s
yDqZYpXvw8qfhpFOqblwX4Dlq1dyDvLkoQQgpQ73NWftRk/nbu6lg+fFJvIao2dsJUgruWyQ/yUJ
4jhEzT50etx6luDkwW4Lb1CXiCvPPyLiMb4LqQL0W5hO0a+zd6HBcOxwUEjjWKqWVgBJ0csMJBy5
mn8XKTG24rXb7lobUO7wb/2d0nFRr0fpKGxkvAZnzePBSMwa2hpLSqbIPPlKl1oP9duUCbfeJFkv
NO3aTZvpD2hxOPSOY52uypKPApn1Lh1eWzzPkc6Dhzkys9DOOtVwrnZoWIvlxEjsoLQ9RqGQItQg
TEv5L+X2qhO3MGcj0H7myhBD6HYfrXF5IEULi4rLRw3IcQOn3c4O4HFhPaigp2s7wM9LFx53xHTC
BvIJRTnRAUYbCRF2G+tRNxjhtohvfC3NZ+eCpQqXENECWGC77J10xNRQ9MEfCoFRkMtXoisz4B1c
P0GtBSKTp4LOK7P4MQ3ta+fYTahu6WDJeBwlMjI0kMmGN9teSc1F7f5CRb1Won5bdjaKwr4CTfBf
ouJgrIooP9EtpS0aUk2rMNYZ5IH7pOH+QfyLmXQCbqpflJZNFOeGsuYlluQKgMvlqf+w37UrHZ0A
fh/A7n2WdaYh/n9hO8OV6IDsOMFL9NHmu68kt4Ap+GMCG09iT07F1zsX7JasxCW5mm/Jgt0cPTnS
2pG8Y7/4GFI7bk0It9pag1DLyWb4RLDOEGQtF6EHEOOrf61r0MuVfFrS49kKklP8T/ErKclzcJ4V
770aQx/sD9CwuSCSom1y0yOdEHVIDaI4Fi5/aFuT2Ac0/fM2yB/ffFo56sm6QZRccg1VKQWcEQOH
DfZgEoz5hj/Hx4XVbdiP35JPBOOc/eJA4ApdfcCzFJV4iebpGX+Y8mkVhDwqolk3qtn1qpIiXFSm
VmlbMG5YFr5rjeXkkATKZ2GzvLTqQzvAIxIzt8klyKiQDJ1PiIloD2gRicTgou+pUjmSKWGmUrxn
2PZvO0CQnOO3Xs+Oj82V56dkc2N5iqeQwnQs5eRGxCIiPp/61RZ6Eq8sqxKfTii6N1r4nCc6SJJq
g2V/2S3vEecw9NoS3IAvgxoKt5Me37Hqz+NoGgYCmoeJpHb/uHnPCqQAuvccJs+2bEWk8yrs5Vdl
04tKj4JKFOB4E0NUL1FRdQLfV+puxspOrAc41Y869UQUnSzUxp7fpQXGTA5zrtjCMqJsy/Kv1FE1
tqLyh8qc5lbhJyahI2AdlpFk8AmbwrY4spGOI4ptqff7Wmt+L5tjBexOoPztKxLFlbLJ+L5JTYsn
YdXUzs06Meb2/w5qenyBDHCyyvW2E3G00yi5xTh72SXs48DJp0gvFzmHsplgJbcw8sbL9Dy5a9P3
WfTNcDFvwQxnkg9qW1e4HTduQRUUeTWIFjDegX/HSrWTfipU5kEs4UfFT5SDwbzho0EsW5MYfqXl
Vq5C1b4RSun+B05gazHOD8KBbPJu+FWBgxlfpsJETu8W1r3wrskcbwb63nYeNnVT218IPbCDb/VB
HcOzaF9mO7bSNPIoftTPRTklb6RBB7DEKX/jp80U2BqDKUdSYFc2/PbzpdhYCb4nwE4G23t28sji
Q+z/V4ecEawN1OyhVa67QpNzXJVhe7nJYfmz031HABTlFTxrbPhIacBOj+Cb1XHPsXvRKrkFv0b5
w2Fj7Ie+uhIYrHXdVK/cis3B4EiDH+M1F3oyfvg2U3YZQHA4JfO69I0nBUKi/WJr9QgnqyFm8hpf
Crc6rmbwdHMg/9qcGMz+MLVoUYZm2eyhaarOvGlFx5cL0sD3/IcPTRWvoicaYCefztpc5SO29xsI
cIp2WtY8S3yHTCo7+R5mN5K4hUWXm7M1+pvoKegULxkvr0R/un94EWqI3NuRFlToNorNpMIIBLZy
/F07GvZqa4fERyBdBY/V/fcWxu+TUwjoOnSlJqCJKB4k7FnZBgNHB79wlwg3X6PBzdtMVJeAicgn
VI2yEkQ9pomxcT5NQc35i14K0doAyVczt8r7A/vjFUBJwIDgVZAF1g6bO881IsqtTUadlnRR/ZeN
vdP9VfBLL/TLlzM9ygLjc8KV4QUSR37SmV603u1R3BBCxWB1hVVCJz2x8BeF+p48g6zAAhnzltkD
4a5Wf2nUlbN+Va+3D6N2lh2LKbFhW9U2CueGngd5sY1bpAryzC9aGAOQUUm4YEgLk5F9k6CUPRoi
mYt6TiizMEsKfiIcUrZaw/cUmbSK8ooPaE5ztFK2OkxcziWMpV2kOkbwncr9tvHwJX+4AthlwxSO
/I51pnNVcSSS3QU5h9OK4MjH0vgwohcH+rlKNspVvLgQ1JF1eVn0ASCawaTwarudMeFQXKEnGW5d
h49CquMlFdQmvv/pVZFI9FutEF/YAExecRGXbNIOC5FiN+chrSoFnkvnllaWobYrvQErFdufbw7y
2oiYgL2eNgv37kgSZzcbfdzlT67bcd4UP+lDkQN68p1FRcvVyHxnqvAWD6z2ZIo63FwskC+2b4Up
yMYH6pcnRMhtzWFnV8tetziXl6uvxJGhVHrYux9XwrJKwcsb8bMB69L0UAxV8nsYsgjcLmzerxos
xo2unxX3WqThRK6tn4PFbuo0AvrJ5Ho5UG7nUf02Ye+fIYIsalkhOkFmC6OZrj4zIbZKII1sLJyu
roZRYNl4fwe9wYFvAUnxIU4/fxgHDGjyBukWO3gUXH66zFDPbAaqSWyQGG0lTCzxEbThV1lz+B7l
m7GSHK3wcmUZ01WTAiaVgzQ64tx/2NaYE9N5TDFfIJ20rNSt0s94NaT/dbyuqem71kN1ewEorrYv
IicsS51h7bHdhY4hA9+PyA9sHJmxYm56p3oQ8fooDiv4qL0+NjzjWydbY50aE/UO6CzIrwZQR3h9
za1PA3Bj3Ps2399ShnXjZGlKrLfby9UT4TH9/U1NGl4Tsu616tiknngV6gV34G1IbnZBUzH2QHyy
hxqDvIZfjmSdGdzhX6b3ONOQc6Hc4UBp+TQoOevn6l/gG3doKEUKnXheYtli8z9kEs8yFN4jtLqj
Gx8xBRLz4C3Cj+fWAZpAWe0ENXKPRKlr5JEC/qyGNY5kaGJbxVbObZPTqMw0Wlh861hq5BgC7RC5
80qwfL/Gy4JMxdL1jfotT1FX4HdLtvxmKvy8b9CeHlOBmsEQFSYx6j29qNoxDFFejlOko8imBfkH
OJGNCOoa0E3E7NUnNI/6RFs5mcKLNVnro0pR9CfkI0/K6rXuffmHQa4S8YmADBBYeoU9GvXIHLNj
NtXcVUNhj7Ijo7VNRMm6tydrHR4yG4JzP0fnyeHrPfVvndTjxUqojGWJ/Elae56ZUHgfzgBq7Lg9
Nr7ApzdIMTlivlS8r7DmFxVgyY10Ito/jSSdQe7UcgHA7c50s1RfYHotVZpBpO8Ocjsfhh1wSTPF
TD2gdrgtxn2CosoShPv/G2lOBDAymn0wzTUN3cWcRYb9DjWk75leyPrruIVV6WcStwrv5xwW/jti
yx2Jw3y8lp9u0cfA2xOFxktVcjisAC9u8oyipvTS99FgsWyzBEEYTpjx1Ggn4JOIhGlAoRG9lCRY
76oRg0J+5CHixVbw2Q3bsDtK362LR13RHM/Uzynign/7evaNiU30IqtUDxrVKAlXp47GACo24bKD
saKUE9S4IBTY3v4RoqGMFsMAd0EACB/es/iZ7ZA7l155WxhouhoUf/B8xhrGV6trM1l8fh3MfRxt
E6PGSNXafIKehuxm8Nju76zwi+axuEBLsnkF5xEA6IjTNluSrz56o1DfKzauPB9OhNnzqdfxmnuq
0woPrRlD01NNIO4FLZkL7STiCqIzWLFGw3vsx+aTqUp4AwJH8owOkFsUKwB+q+K7fvakHa92KVuw
w1zYeG4TEsc6r/KQ6dSJhhL4ZsFo18YiN1yOhxy1duzqSeaFpDNTWSMVZKUUUiJ8vLiySw4mmn9s
0TwOmQOw+7TXojBJ3sH3z9jMdVf6VbQcK5xOWmuRjxqIPxxHsrkrYDvgtydIA2Ny+hFx1/zeydU0
YQOhe5QfSH12lUdP0kHhj03Bc4j6+EvOF11CwAie/ysJAc/Y4w/mk/u9oAoGuGKRLSKzsNAWDj+f
HSlZXTEGQrgkwQ6YzPWqZP4gCh3KVjMKu+JwX0H9MBrchWPzk4syX+CvvDkJIpPDYvvFl3xgPn2I
+Wp9/Cf4/bsZt9tieoIkkDP0JRZ2NPyQr3jNey8k5WLyJl8p15x4Jwqql6mX/Z6F5FFekVbuzJ2/
kt52NPr4mQONec95dUdcLUdanZYXIWF9ppcbg/s0n/9PAsVn2BE0D5VJnASmz8dWgr2wuD1ZGYtS
FSmiSSZwDgNWv0ZbNeyyySeIi4n2GzuO/q9WSRClQIEROwzYPl5AhXmkEaVInzj1wLb+7pnpUxhi
Zs4rdo7fEFIV9/+r8aSoJRgDXkmAifkeYzhwSdTq6yf20ItOrwyuVmByeSThA2Qw5kX5Z9qU9gZ/
4XsRMXjC7CdmLjKXr69JUrprltObDulsmshWCMAy246D5zOie0eTM3tz0YJ3xWNOwW7W6rXFknV+
v/EsG2Ne+paFx2bskQHJddrGXVCh7dwZ9CK5dcU/z52cjenhHqQ7FdD2+dRKGZ02cr1LGhTGT2rQ
PUd2j12yusRwtJdbvh+0ZNpcLR/zUEEcLtAOa9wVDFeup+5lmo0XdoOOs4K2tgB5rELcYeFZJ01y
ppTdHVUpNgnHsYWngVflTWPmqACfhWC9omt0kO3Ie/mq9GuArI9Vgamxu3i0nlyu6CuiTjb1rvw+
Ub2rEwWVIDhz5P2yKaPc3EAc9skH7/4CsQJatmPBfR97ZkomyuLEiB01CSe3+mKOLm90/Z8l63YY
qfWJ00PWDe+twqgglIBl3NZLRXM+JevJgnpY2WGy9Df0gWeuxwHS5Le14kWPziTPu/jfbSBvDi0Y
jmNL9aWQGumi/stRw8hYrPNP/dNrtoPgjaOggFMXHg+mdWVeCDMMkt6lxRNgJVrBZzkqxHLM/uc1
TtAb9Ey3tOF+tepn+56g6rdEofFYIhAts/ue/BpBaoeloXkrG03nzIIR7TDzawVX213ZxYKdQ0Ff
Gig74yzTe7vFxLEb2LhCs0C0asGbjk8/7c1h607TaCdOV8uLBwXz0mpYVTGOJqKYcTrroz6irChL
hb6YFO8vaIVY8H2symRqWgSywx4iYETMnR8XGLqsqjOX8gwbAbQ2pvUcKcKTa/35OM6vwoVuWhT6
ygee38BdVARA1i/T0K8dnUOIJFW2ixEv7sDROglx5DhZek6Lv9G06JpQ1YEX0b9XjdfIIZDZbQLq
c7ij0Jh6BI2t0SjTAv9XHTH5xIMD9ziMezBuKMD9aVOQ9/JJ/2lm5w3WTw82Fktnxs3Efl7TGQI5
rftIy7RT2K/n/KhJpLLTUfxte3F8E3vGZASL53s4bnxyQEqgBq0bWfcYMYYcdaeS+fGVs65xDwtR
e4pw2qAqhlrvzc+YdIGyYsq3sQDjT7ExBumRQPsj72/MnWbTSsQfJnr3JDN1UH2AB4+2odbsq8A7
iX/bPP9CbfIq41WsP2gHbBYzjsW6ViVeIb6nU4L2K5u1KS9ySqR3iNeTAThJKSIyzPKpogB5Zsg3
+sKccsQ3jEQwgfvLlUpl/vklYo7ZjV7CbcJlKufLzYmOYXunkLiLdA3YXpy8VWR+g3rcGMjI728M
XdZ9DIhOn45gNOa0zVCdBIrEV1JcNxfbU+MXUAyPbRlkyQIBqWwGMozpmHPqJ4kSsIJo0WwoIwY5
ekeqm62etGnp1V7PE9e3ZtQIv6ta5EW5kge1pOkr1O6cY9V/o9TyXZozYmyi+IS8LAoz4f2qo+gq
JP+uYfTliY38j03l0joUKXWnvkZ+bUwkx4NZTBjawEYIxLN0N0lAozE2KySIHMJNcRivh07Kp4Yz
xh9nDvT+2xQqxcOFwi6WQ/d+Tx5Ge6P2mhbqEAZHb2vVzep2Pc32+SlN6DDq/7xXaNi6RYILg8qk
QOUmlKUy3hX5fzI4EmUmzaPqif+kuCcBsiSRQtIcJR0cgzikrgsrgcTWRGvb4huYx3Se0vPd1xAr
w8HZ6yupu4/2zuQo1HIlBG/u4R3rFhLil7y9sZJ1FFhS+7rgqTtlsh4NGsZYAc6WTvh/WD0FVTzj
oF0FyAMmK5CTlj+hkxP2WGu9W/ezG3tIoAiFRntvdX/NLKbHqDE+Q2sINyMcNXgOGBwh4Ssd+2z7
t+u0lrW1WLysB08961UHim+xqfSdVZ4CYl+wL6n7n/DHybcKPqLQlVH8Vy5SVNMNhlNJ6j/zXx3b
zAU2SCSMJSBm9oSLddxQEtHlj3f40sU2ygrhgx3NSteX5y7Y+AkNPGTbPW9t6PobJxarTr/2v+M3
p1gdFcsHO7DZmy/GnFyBKTmWXfUzLQadmFW7BURRxg89qMW0KDZ6fCqPlM/3KZzl9+vqVcfiFZTx
0BUkhAWHIIwDjKDYlVWXHLYkrFOUJy7W3dDLZXXg442PEjA+OJC4oImNM3s0OyX7FRLKwPIfWeLx
4gzxb9Zsh+UdpVJ72mw3ZKxYeqLDISkCfuLdMdFSD6x/zD29TcFcuWpL6tv4l2/m9ljhBdL4odZN
kWRO/xaQ9YfXSy9y19wYJyDalAFGe7MditBI2ZtywaZyTpzhK0CX7Fmfcd/SjUnrnlXsUc8FtH+a
HmhCdiBwDRvY5jIVNwj4aE81tfAldoIY5t87tJVnZt9Kuw+a3ltYLS09J4eMQF4pt2qsDvtwx577
FvnxL02Em1k78JdW8xntd8eW7pcEkaGVfiXk5Us/iw39vPkn5FTr+0Ue/xvjPBc7Sg0B1QOmnI0V
d3oX6vIwGRab9M3ZZbvW3rLF6cj7pSLh/sAg3w1ZuZWZhapHpfJ52qZae2thj1fhuQ1shf0WGYsD
1GyDawf6OAXZz/WJwvsyCYucqDxY6H1nQourxcE7cN0xMJLMCNE6RLFrE89bFFtTupWsSeisFn+Y
+1fu8iZwk0YLqiPOL4HV9r+mbK6sb3fXnO35Tqqi1l13CWydOloM5trtrJSvuVWOjhertPFacm7E
b3xXi3RWIg+XcPLJvkSRtL16e9Zi6MMIBP5ZnQYUPS9rlK8ThGwZvyGPQwF59I+Cq4P3hMtkZ2cH
ZsfiW19NGiSOfP56al8hVP4Zn8sBPhIgvlCbfgFOBf1/m0P5RJEFwSyodLWze7sG3d7b1Jey6yJQ
1hf7NjLsjtug9y773t8UQkmOJ0ywrn7BY1WxMT5nSbJsLImwiqApXdF+B6yXJERduK+OrdXZRZz1
ToYmPYLKydZume5bUFr/dxEeG3Hx7MwsvVeY47HBtpv4HlAUWnOjvD34W+DlnSKomowLdly38uGC
IF8iIDSWfB2iA5e+GAoeEL3SGEmFXHtGf9bbK9xT1N+xDLKXRlLwD2+d84YAB7pdRYV/6Pqdlz6O
V703vbv0RWJymC7831q67qoP8VXsAF+FaCFegIEgGcqYEZ773iSKHT/yKHPXp2gu1oWTvpP1bzZe
k+gh0T70mQVh1H5ASYvvgZCmGV0Poa6Ymwdocjbef/dHF6O5NMDLlrlTkePVLxFT25ee9w4A9acr
nJWNFvA7KqLRR4vjwR9XOSdRiEnoHs1GMuhUOpcK/hSYvnMJ6rktvx0COpe3Dol9Hw6vEnVzG/WK
mnQ6eDKXCd0zj0rOjzeBBln6U6lVbW2H8NISSMmywuN5IBCGq6ty6Ri3+EVfuA6F02x4xOh6EMnJ
+3jLj4jsNnFoWGchmqtr+s1VpS7UPeRBsGGetrU1ic7kg/g4I96nhUs+vM/8Kx/gCtE1O3qdWe6G
tcplHxqsRabReqiqg2DKVyY9PU4iORLt72mUbSv8Ayyk6xKrYtWaeUkWDpEbHXQqv977bOqBhkny
Os54pHDs0HDOYTGEN18W8sRaCff0xXwHsOlXUtM7mIVmuK1no/q0FQUTL8AmFUPnGbzmIRZ7zyrO
hz/HPdmKIhSADNF++bb9aSCxwrPw3nLDdedQojQX4CGaIbbHMvQpf5MWxQpru7GtCUPTCwBLqMG2
dlgHe/y/U1yiQz9RoVyOd3yNk8AbhPcpNoK9+cchVGhMnY1Q4Xd4AWXefkQ/QXSH3KvsWmkDJGET
9QV3VaEaxNCd2MzNNDoHCAwliGETPfJPlFQ+1BukqpHQYNrDdLI7hXcjZvvELLkcasISVFgcnXzz
KEf2bonOEKWIK5qWk8V8jCORa25gLpEgAu1cpPakf/KIpFFhrm4L/m2dpXwEAHbcQ6pvsALiBFf5
Hx+UhD0/aontvFo7ERU3a5YhH9mJvOfjKq5eindWd3vWm32pGapNY3vTkhCfkT6uKSUdG7zF6ksL
bMAbLuVhviOiwZYszbdeK4s0O2JOmK1F83kJVzQQXcqLxNoADdyFc+xom/P0an6llB+KWHC1oNEK
8XPyUMjJYwVT9u8KnO/F153RzHiPxPHnYEXAm5LCWw3gHhKSMth73NUw6hpBLqTOB5ra33fpOtwb
iKmpUd3FYLPciELFGo74GtYg34CVhTPmC9s20rU+HHiuSoXu8iqNI776dba15dQvwg/uD47SzUmJ
IrW8bGs5IR+tRiAGvgcZVJ95UlZLGEEWHWUhVl46YGmAwJYlRsFwKvSqCVE2w3nuM26VivFx9pUh
VA1kUnGGhEys8WhDT4fdSEC9201jgRnLZH0CtPRjpTPT283Pcvlbhn4XcoGdulGkxr3cHiI18FSL
Uk0ey7YPXasJxmf1JUyubdvT6HNp4tVqd9kSYIuDlXHTv1LCkvq8FJyH9TW94TI55i9R/w/Xnkkl
UFobi/l+iYwY0FDUUFOBPqM4i7aZQ2CwETpenjTX4hNfJ4bAhwHJMsR35kvt8OATk5L1SnCPk+Qe
skBzjitKQqCgoNCHDUThlCtKNLaGFuwaWJQgDPI2DwmcWQT5Xq68LY9VOZBPiwKNHM1fEQ2xDM6i
0VEZx5peH48BwrpKUEeXhCAFE/BvPpvRFVCxnFpu4CM/pW3wud+legurJ/NWw70f4+Upu8SJmRiF
Fk0IGubOTNRpvfbNzy3k3QsxrsBRp3on8uyrkME9VMDy23tRaWXuiDNyArGtJ4PC7daDKkOouBL6
cahTtfZOoit4kO9jAhWKgndC+jlAB6bXfWp/PywOb/EUlDzOLaw/D8vmXUjOTRittui5u1QUlDg1
jP0FA1VtTKpIDLf7m73GU8rmjpxLZxZlI7Sas4LKOQN6U2udNsNZm8TWvlnypsvhWKf+zeot56di
7HU7s1l7YVNdAnSQ5XNIUBoenTAeHzeeEQoPtwD0D/7cJ85heJyXyyplw189HJZDYvhb8ilJUWwk
Id3OSiLrGFr8U6IfWO82xL3zg8rNDvyktdtWbkiRONyiMrKq03hiix69kxQ6JIJqkIFtEStaXvYR
L8UJ+xELADIk4vnJ8WaVTqgis/1SJ1fIRM0WJK7nWNwJJsOdmOovj0UohiDcZbov4SSxkG/AzamX
56VXqAJmVQ0K8uOQ+BfMFCWp2NoXxRS4NNleQVIFVybySixpDCNc18ExiCTAEzOyqnls9MM8Zypg
K5EZsICRf5K8VSd5rnt4sJeucpLLjgyia9LWcj/cZcg5oa45ha+tvvFoRWp7mRDGSfeokfp3SIh9
EZZ/xov4GW/3Elly6s7Xym4B02VIpntImEPbvYM/kH5cwsTCgblPWjfe7Lc8vbJRnI4FQKW5EZW/
O66s4gRsyB/Wh5YMuKqpbozQhUAirayFV0+tYnuWIsUR62x2g/LEBRORum2xLRJAUPMKZnsi9A1T
dsn2bXtxYOrLRkhS2g8nXzERP/Vs4Snm1DeRrPtmZUGs1xz0kpH6S5b5HosND0IMmbSIBhFcjy4u
dJnotsJ1mWrMG4wjPMm33KD1cUitr282uGBmrNAUDeVEsZOxHz/6HLstVqZIc+xSp1yOL2CeLtfz
vfItjGCA+ZGSvVJKQX92rTxszxcUyLUmwXgGVi5Tdmlsiu7W+3gZkbOT9KgxVdpiHfmlrI2vfVkt
OZG1EphrxUSlpysBIezICOhUTxfK3jCS7sqiR8rUeHpJcuiYHCP6vMM3z7s8iR8rsmPnAimkORp8
9+N452oeVrP0LR3dREsASKSl4pdrEQjL12Dhmw59r6l1y8zJN4aIm2ToG0WcbRJd4XVSCSHw6/bX
vQAV5q+0uGwAhk0LTXYfQo9/MsuDwz3q5jxsEf8NBKQ8rxRaD3G/l+KAT8J0tDvRCPDHKSULWMhU
J7UELe6hTFwuurewZMpjV9PapqpCzHTxD4jnySHr4cws8779ok8wnR1vhGWy+LSOiQ++jQ8oojWl
uwXZ3boVKneYZtxSV8JGWCY+QFoFCtihyV/8n0GSVii5UFWNakpxkLy3El1q0sktYAPCIJDgNcGV
xaHM2h/UnQ2oS7gbstNkeMxHDRGVpS29gAVdC8qorLulsoKUX9Dv6odJ2RdjwYJk2rV2cXttkL8m
zhueu2RxeaE9y2Z42EL0S0IKIaytHIPFHi89DZ9WAaTeGMlVrtN+8+F5tBbvYURsluNhjrYqxuw4
E2qiRbmjAvkJpist3wi14QVAZkprzwDAe+OYd1LHXbO9qR4ysd+mk4AJ0pwdKsIzabf0q9BXVGuW
I71bONAXk60S8spv1A441IWgLjtflONUVaHql/6SUzrVfL3wNTU9P3RCbLziHrs8ZTnNihtib0GP
955olW2yQefbiiS6+S31aTnX+bPWV0b7DLiivKtsAiEMVkxfClDyE+qeq4zbhy0Ay0K4B63zEpJ4
cUkC7DLJ8oERdqpGOdomAhkCP4aXuJGGWgVS8nNPA3pNFZoKFB8RQD9ive9AVrL3/QA6Yyz4dTWy
c3iNw4S7GCxDe69Ls+1YtBnrwAKr/Cpe01ZQ3J1yx6YZDG68M9OFrwH6aFP0wKm0Oa0ljrtB/fdx
Hf66fj/AwNk2X6C6HeJTAfpOwZk6m0Af6sc5oT6ygJT3F58aZLv7YtMwLGv1Vffk6aoCVVEkM0Aq
OrlNG/vXcSGD1p7KHbW2RT3TkecpmUZD8xrHe2wP4uypahNEyWyE8I0KjCCY3mJ2gN4V9aAm4n/0
kJ2rO4ximt/EyvgCj6B/5dZOgSYhye2xs8D2LpqfYJreL9jaYiYvYfDNtrwfoS0iUXc+Of7gb0FX
1ktdWekXKsEvTrw68n7kuodd/NWWPDwrnoBcRJhr2jFFfw1hxs3GO6v1LVvhBXJX5MSS9cJelkCu
O/N/oAVQehtaPLkpwT8591sgThcLn3ulmiBcq9W3Sff87+pvPwxOkK3qT5Kp3gcfyaKIdLap6dKG
HkvYocCmKJDpRlauwHGagcSyPDzPXfIrva8vFxfXxBI4zcmD9D9Rb+QiIBJAiplZJmukLZ9/70lD
oClaPySBEC7+EPe7REwwCt8P1eWKsObnx96rW4AUUQFO9noqGa/c8rBymxOC0sj6LaQl2xfAyb1w
0EgExOTv/1w9H6Tt5ApAuCPOZqHjjXw5oOjCtEfghRihjmlN8lY22xloyklQ6Njzd3c8y38kAU2k
QBRnm4PaWeJUkMeveBzGjkN5NZ+qaujzDVNmwYJU3zvcWhEOXsISWHglZLlMR30xgO6Hw51lNMgJ
yj5dKH1c2ZBCDP1KyZrcA/kWGtFgGhxXfRzNRlDM1SR2bR0mQh64so1zBdg/ORZd0ufQAv7ALcrW
uYe1qH0Px8sda+dAA0CZ1f3Kl/0tB4kEnlGWSEiRd9JpyyKp11IjdvAeXzfmNdzw6n2AWISL1AHZ
I5xd9JyAyxGbZdr/c/A0zakqvhyv6St7D4rqHwiyE6h7cW9VohsXwUY26L/SEe0mpCbrLMAdJF7M
kWiM0JlnilvqYoWGbC80Mqaiko9Q0XgdKPHb4lsJNS1S4DsQnJ3DWMcqcaa1kJrOql5V59SGTJED
T5TNTuchGnDpCuSWpYOdR4FdgFt2cuoN6BtAQHuSLpIcnbdyTuRhIlt/o+T2t5n3VhrOm/3y+xNa
wUSv1KCCoI3qrT5MtH3Vzpah3h32vhOiJZEC/9dWlF/Y5SNsnP99Y8WutELG5pAE3jYpa1lXG25n
VBTiOoD484z/+n4qCu3YBYL03QE9usS5e76pnkInoyOuQ6ftzep6hF5uDJGcthqTzJkuG9l64VEV
XQCxpji5DBXFJ0kmMRnRSw5FgI9+kDfl1czeFCmvpi5n3KUbIKiY7e11IsA/dD/QO7ecmMs/ChAy
E1HYmhd1Z1DznSVgdJ+MmRYEPc3FYZZafkuKR4T7/n89AlkjqE3Couovh9l5kV+3g0LJBXcsuM6d
G0D8DgDD4Vc0ODesRUb0JkrdqEWnzTZDkB5CjzhnPAq9L3a8wYSIshJ1vmUnsjcciW5bKL74Vod9
eqo8xjK26+J4FeP5fBb54kLTkXqNyuD/kymfJntsa77ZhDH0oW5MdnypqIubeVMSE3pd0RFvET7v
T2s6SPD71M3T0BlCY2zFap1lwzLXDy6HIf3VtmNmg3AzP/RHZMrI2M83MO3YUBStkPQ21Zvt3ZaY
9eeAO+QmbJCgNBjY2YLAzuZGz2LpqSp4uTuuNSuuxDQSa9maM5xA2pPfbUkLmZwhfDoGZwulkLcL
H2m09dMnWQKI+iThyLcI7QkONqQcrFV0AFxJjJOWAM1qVkiGSoCfn+et3E1zX27Uksfvc32uQ07I
0i0DwgC7q6B3fkfIjkW+WPYihg+qLJs/LBK16vqihznNuClllMvJk7kzGfBxXBG8WywYzKeigeem
AgAWXvftSRekCYtjpmZtw4UTH7aiGYrvFvpmA561q8Y/P7R69XsQdXEDnQVco4a3+d3hg6UHe7R7
+jwC1xXLXoXBQ9jd6b4Yp0zS0ysPn75T6XRhR8d1uLlVhbn4MxxNOUzqWhtVmnJEt+1T8J2afGUh
0J1klyyY7u+a9AtMYbT6tlk74yl0vQmsmcRYbmvPDaG+qk/j1AH40Ihq0m66EEoC0YKERjCFz/VC
lsmS9aQ2SmeLx6eZFgkguPwlbPoFN4RB/OBgH3OW65/agKuTItW4wvWhj5aKwo/cFblghtiUckgW
9pBqqP8viW15CLovgxc1a0abv8/O9d5+uxo4rvOo5slZDt92nCBEQDWcuTeeCltqQp63bGbKQx70
tt7g0ONoygoDyVwPlyF2TvsBuD0Tf+bCx1y3jHKr9k49FzWCVqJMjHCSQobXp2QjH2KLQg+FP5lr
wDP3I8rrtx09U9zYzHtnA6LI2a63vWsncWpcP2wQMH3NysZwe/5v4BYLcRfovnF0ysXdF4/uCvi6
O4JAkyXaYLn/b9DkjFT9aOEjI1gfw5hH+hCaWFP0knAujvoqSm2Gw8f16e3p4CjTFGD/0tWrEcBZ
lR8wf7rEp9SCeRnSKB3MrkwtfobvUGR36Lnv2HfO9KOiaic7/4krnV7kmEDmmSAeUwPsgDDlXFRA
D9XHG6N/PF95QQhWPgphvlSHm5baSummazcr6goGMvrmfHrmXmew9N0cCFmv+H3anwZ65W3F3OnT
MWQevDn6Lba40fa201fp3ELGyohk2kfkz4tr7xLmc3dk49Vo+azObk/xHjQBFLGnzbXKz8VjIJ1y
VwLMhJM7QsoKNwVTrlQtYyt+Y4n6dWMt1gaxSp0tHXcIKf9yyLl+T8TnJ1lPCOVyeXx3m0Vdac0S
jpDInEoTY3+nGg1vd+lAfr53OiZA8tE+AbtFSu+jEpoXoZZzNmoehb7lSEwESDlnJ/7zZFxoxl8Y
fbONMPrATfrgiaPznEN0t/aORUJpwTRCpvMlC34QSxSiB5FGOMYMiXX69WB0bbiFBKBWd9GadQTy
ZSwEhBnqnsr68MtSBNZiOwPhNsKkwm8rWve2EzObVZyC4ThVuFPxR+1qlRu/ax5so4oSUPMMJgeK
vLCRF1iI/y3GmRac4VCvkOm1mUiCdyS0eKUTYbQ4lwsigrNwFvSsBzPpLfonTPLW+HioaGhBGIJf
HQgISfNpvQT20Kv60PeziX7cl3fWau+pg+++1kuA7SncnueUKYDuf+jwT0ZuqQwNs1gWb1pGkN2D
DBYwkqa2x4YMGACMh8liUI2DUsdfYKYkMJhZvIVjA5q5wn31kIkWnQxDBtNUQ8LpRkthks/ZaYjn
IEzj2WaLBKSNNTUlONnMJ1DfHJMwH7+TNXU2IA7q1RKmQP3kWvdiIK6mC82SpTCLdSAO/73x3RCU
zPqpEqBhnyXGyi2LLcRHImfoUoR6bR+ilTrt7S7o2/ZlNbcaomGFOiWIrCLOrfkF5IdpLYA60saH
ameVt5YgOa1hLN3SfT6GBGHLxFEwzvTrJZHF2ckQgX/kVtTlRdSEFX7MCRCOXYjUHa/Omx+eW6d9
1nzQD1g+QSlzi0AtVSGTfeeB14ewYFuLO1ScLo4Bc3aOVtkNLih8TJsRt0ZFQFnPmraCO2YMr+XF
3xQQzjayCAOf0bCL1pS8fjQyUXWTYA/YiM881HDNx//jELXYmbuuR4+Lz/xCL6DUOMqXMPDX9MyJ
JIMSRtiRS9xpCzMibAtPP08PGnam0vgy9bD7Gw+e8L+MpZOVUS4y4Ebgh3dEzuIdUL4/SPm84I/v
pgG/kavDO//XaeHE/fvrBxSVQ0B9JcoKk6Ir0Xt3JULm7fa+08xGvKdX/7LquezCbLNjiQtVczfA
dhBcrQu3bvhuEMolJy6pGD0hoqKBYUJHsHTZPk7mryJPTMqM4GJ3XNIViygb2vX40XF0BA+Y1qsO
SMQxPUVfANoBtYr60lKsIh1rqWbLYpQ6y9uqXDcERqtAhrJG1RjfWFVOxV8BlQxWW2F1d6/z+2/G
f+swMnYYgn8Q2vtL0pWIeDouENLP65VVg4mjzJM+Mn09DXWy6bmdnn/LTqGXHHJPunmsIcWSrdU+
Zct2X+NpWaFoyyKNnAgPGw8HQ++sFv7+BJWXfBW2AAH5c355O/vq9dxHIlIXsHl7eqFoISWd9OjB
DJFqFDWzkUFgAHVuWaSkVseInTZPbHRtbs/tkY7777wwtjEawE+/HxL4YsWL4rCYi2PwsKYVGavH
P2WGfaCFlODdxl9rK7NAJRSJcmV2dmA7RByO5Xw4xl0lIw2VNSA3ZtQvOOEmaqnCOjrtZxdK9P6F
xIG1Tf6kg9Dzw8gqqYss+gDH9WmKrVp08eO//fLIgkFy6OTNtZi1zyyg4rhYAHkNNykb2tbZFFto
oVBuMFDTsZ2DtnJBX6AcneoCN2RKTMXYVaBKcaTEbDT8PLN+ViUIZB+UeoDU567xqIjd3cnv7seF
XSLW58NtEvLD5bY0n+lLS1FMyZVHXK4Vqi8ftLPQ5SH6PhztTDHPBGVH8vYpwL1cCXDi2eexSG4b
o3FbFU54tcj06cl117jeLGTjX0mcfpGIpGhVAwyoY7rWIBG8Ty43Z1rS7SeFCXgEBQBKVsWy4N3V
ZLPd39kO/h1nv5xwLeZ+H7KotKcNHMaHBmU0kvQ1Da8OCeLH8KeKXxYVQtD5Z4VO9OnbSujblVkf
ck/b3YoezvOUtOLudqiAVZN1tBseK6M6SLbfKLoZpzlWMGfOB3aXOUCzDxatLVoIzbc4+m+xGA1e
ft2JlLMPfLeyB5XUEird+qmavudIEPNYUz6Wr+K4jhqwZdeBFnCl4l6a9fBUJ+0Zo7yrTxF/6zSt
b3M+IwJVEfbdVvlqlDZqhDS0pc+1jqyaIzdKxwQ2Qvjkipj3lN+2Jmuruo+2liCxImCO4sQOYNyy
/OJ3XamIqlQ+nXu4mX8QUgeCKQeFOyIDMoPusRxy4Ti6OIZtRfzofG3C5QuaoNifq+Lhq82dyeeE
dDoMQJHaKvK5eLo0sV+dFeDXQYhe5JQqmgbkbqctQscg4c17StEogt0KO+FobcmEMqTj7dPAFlN7
462Ic/RzGb5Y50J8DECcCgxwakmI0bQ9RMfw5QIttH9ZRyCY6YNknSoxbFevWHndlhKsyDuM2CIu
dF7XA70TcRE1IlqQeE5ZWYd0XBkkYEwF0E7bzT0iJeezp3R+cXQKxmI1CRQ5zsR1YCzW3XX7f5YT
hQz4JpfqSdDCU99YA/6jJ5zKH3N1bTvRV3DHrJDiLNtnVgm4dHo5P/S8tn/VZKm7dzeScxn5fmh5
dzT7sz8581QIX9g2GoroQp1Zl8zo/MoV6ycC4JtKZmeCRNLw25AbdvRhsdeNnRYE3aI/jNoabLbR
7A8HptWJzxPsdbt9tM1dyOe+Sp17Ood9lNWrc+dilxQp6oMDnhAmfx2e9RKjgAOfZbbvUNDYzWad
vjyecY4vIYO2YHLSwMEoKgbAEgpCqU9/u4R9z4QB3dpwYWv/VeBH0LTgrmQlzLq8h5pLeZGF0oh3
5XgjbZE0+oSz0C82mb3wSsP7CwsBFJA1iwKHizz7T2o/G2Dp/Wtt5xib31V2PpEI5KzJo0uK+jsN
vYHz4uFZ5LrWLa57iVgxyfwSi3L0u+QSaVdc3GYNeyMHuvpU7xvCMK16NqS5tmko0ZfBQJviwBuq
dsncMX85fCR8lY2bTSwoGdGiRemp9mSE42OlpsKMdBXeGdD1vWVacvWw1Ch88muglvfThJVFfdzI
IDSmX+B0N6jX+D6T1NGWZvTfN9h+B6mL5eT4KY72SwuhroaW/koakiCu0G+Gn+RBlhZ6XzYlLzFa
Tkz1CoFa7d4hPgckSZmQPZLg3hNiXlRhryC28tjhIVsBImr/biJEueQy+W1TdZ6JH2WE3wPddc57
MSdyXXp+1llMPsTJcH7Cyqg/xguaCJesYYnKGR2LG992FpAijSneA5AvcPOLInwBXWoAszESkgKR
eBLmc+oJDEqHiNMBudyzb15yA3nls6lQHlWCos0JgR/BnGt6qLNdwjwYNPJHy6mSeiOk8uHlTlQ4
bFXxayrl98x4opacmiDF7+dhvpzGuFXU+OKVHEBMCMECHn+ybAuHvMpWz3ocu8DGRlDeG8qK7py3
oDjsUF61s59zbIOic+qEOJlp6EZ4NxCKMrYVIy3bhZExcRKjVZOZzdxoDjQZ6JnZNKBB+y7pIvVE
c4dGlZHAOa3jI8tUoPlN+vwmFkB9/mpFllIA9g6/duedg0b7lTwlOXhQoInqtA+fxpH6vBzAm2Ok
i73+mBOPSc3UhB2I1k5skuaxoZ/Yd452L3Z9S0qbtQEk/RJ+OFI1dZGKgtlhwB0Jn+R51HKGjoYj
Fm/r/2NJYBIaBqVIXQxfiI7CoeCK5xXAJJPWcr9bT6oRN7LTlYXrRLrSWBtnieOphxDK+mf/rVxF
Tpr2DQXe/TtzBJPA+c+4nDodNlOYPgvaM8UvZPG5pBmKgkao7QaEyboHMlOvIlCNMv6LH+y0kYWL
/R3l4WPZfvsUpUutMvoqJiFPPUxZ7eybyWbw4JPvVG5vIGtPuY/ObJAU25ZwRE7AtXMvTNsQNShY
C4jHK+S5DZh09thEx+2GxhGSnqKj3W5rLWBHeFscWXiIZusL0o68TYIFwS85yTeZLI7tlBYrVstk
KlMzrx7Wb4xQe26np+4Ki7UXd2mGzC75NRVjGoW9PFQGBn/q5s7AY7lDlOSuGblQ72bVVWHrTOn+
SUw0DFmaruSpf5ui/r2Na0sfI6jySZsUI41nGEhceGYBL6XeEIe+jBHPJhtVbm5/iFWknc9c0Ape
Q3PToX4wDeVVyVGdlWNIkd7psDNm4d1USnn9GbaPV9a1JCftTqXWAj2J79fmCz7TfaovKJzBnj8k
M9Oks96xpYg6XnENMtPzaBdG1raAY9QaNPYhoUDPRSXy2TV2LZtukqycagXonQ5gILaj38fIuXgv
WKYYQhVOIiInpIg8vH3dIary0Ivfgw/u2s5USxG9JyiT8mZAUBIFLrflzjCkvZKP5s3Zavh87AyI
r3XKRtYMkRn/RNBb1kZtUCvWzf2navrZ+irJOf7R2U+gc4NVFgPbp55dLkKsBxuwVzN6bfIA7cQy
M9pulm6OOzHIQAUSmNKgf5k/fd2AO/CvygmDUgVqGgP8pCnqtcV61qXGbA4nQIJC0pumOKm5Ojgw
iqBWP81TXJCPVXFOlfqslhaJB6R6uAy7IpgGiFonDNLAjwbN0qZhGbT2rGlZwAzI4BTcudqhoERu
Mi7aeUwC3b/JG5s452fNzkJ5lX3IEUKMlLTAWs1qZ9t2hI1mvEmp4JrK2p8pyil9XSjcicJsdTjJ
YKVJUyhTEtTfliID+FOeppH7lfatqvyfpDl4tOxc0cHdDWqof+7LWpUW6PCyvBNnmL07e93bYvSj
PY5kKhfe9sC0i6dnqmKmrPkFd7YvEo1UoJNodRRvAx1Ple03VgNw2gkYQ/bZw8bkMnwuXu7GXtU+
Xa7JRjDxeMhhHuF8QL92pHcFmwByu+ZEMyFyKH2HYSel/15kBQ8iDboXSReylu2CdM+RCsMB7tXc
pE2DAuCALa91p90iSxZ7lON4iaoft7nfoq428O2yOVusmzzeLgGjAsx6eA/BrliCaJSPsoQiPA6i
7rATDFWcSaZg2hBl6b/N6YNSM8ZF9L5zPL2B9cW5t2dhH/wFu3tI9vs7tMotVlvplQ6UrSvDB4mL
mh5ixkTHrYTuMpO7gEhmuNqIh/ffDI6K4peBj/+lQpuCah7fxdsroc0/IVc3XGfrQFS9lDwPphqz
THeUWRClGXFT9oDhmNZOsAokgcl03S6Cmh7RR0KzSz3DPTrfC2WBL9xwKO7JFPZKjBxfgjtbU9W8
/HmqsItonmLfTlM4+HY9UrhcHOVEIFzJ88E5AMnpb69753BCBgZ/HLQNlk6UCAvCUvPCmdy9UAcY
c7HDBZNzEzVGGSOtejoI3k4uPK5xRsbQGkuMkExFPoR//RFSQVr2IiJoGff29iFMvr3ckTUnDdrW
NCsS6RYrb9piEnSxab6zUYFa1WoKb9iScA9hCbBE1hvWtLogagg0lagqfXhONXWlMnQJqEP1fKQT
iSWFP2X69JiQTg9Pm4xSs2Ecv8vLMjM2GXiHSqnd2b6GqZqDfPWOpcZ9p5GwVQAo9x2vgtWYVn9E
1jeoeWvkDknsVRH6gZcgW11zn1sn5xF9KGMFFiQggu/udstef/FV+/UU79yFysF0wALPr1Xn5YRo
L0lbDQBeYSU5YqrH//s0p54ds+YCMxIh5iCr5bFbwQnlqvf7ny1BXWeP4N89VkaSUVy7GSHESvXw
OmdSojX/UCcMGKdHmG/A0sl7n2t/JAfWaElc+iG/8Gd6bpBfo0dhAQbPy1BFOdS5cfc9hkOSWgNL
5Spxakjd/3KslstFUvkaOh7oyEXcOr8s8EUPzNR0MJopUwS88tKMDb0alC/Vq/kwsJMLU2QKB4Ya
1HTCS1fskbffGCZT+r/sMFbWAbFsd/1uKQJC7xeaSsN6XOqd/E7fU1WKXSXAs+SXdQpw8pUvZK5f
YpWBOoLKRbYfylAUAQ5aC2RSTKYJoUb6F4qwddDiY1fReFLSpamFb3p0F7XPOJQRpA+xODaLVXvh
koAUL9JtErjyeDyuLBkBf/tcSJzPHnE/ev/QstI5xAHOWBlQDOpC73Ag9D4BezCY2ha6xwPSIizV
FrIVJVgJ50ediYxwI9N9p0HDPcIrLsxpdExTdHx/l3jQc4RgCw7B3JKu9xdbk2+tpNvTkEXiXr0e
YE48A34eaEDQstO+PVML9GBXOamEd+3nEXD1DSVe5K68WF3mM1U/rZyC6/REuXiv347aCXy9CtEY
zJgpeFWHFgtgJjHvlHdY+SVZBmfM1GyBn8BULXwi/lyhEFv7soJaG3A+lvJXMvRwKeua8sjJaAWs
uVJzTnkWcbN91faq5JSLqHGaj2EOcPgeZ/QxH7dqyTnhE1k4/23Ex+RH6GfKbWKK1nHHg34C9TOb
M5t5RpNjBVxeJEWknDbVsdKLu1Mf2O3CHPUnLqSjQisQxDE+HB5ryY2V8/92yOt0rwatPvIJ8SV4
cdr42/fHZL0wVogxxZuFftAMBWvEjFpv+OA0pWvkxZ+GWxCczcA/E9+DDGqx+xW41k4KorwxueFS
rA/GhBhAMM8apqFoSFRbMBiY2EM/0nMHAjsZo4ruhaSF8yuP1wetNosMtSAi9KwBJCdpuC5KsE2l
ico5IUs6ks1OFVWq75UfYk6yigZ23I7KsN7Mr+Qns59LsDYlvmgdA+uTgNMLQ3oTcoscclQvNSeD
gkqOsoKCJ8hpdQcj9EACdMaPzrOlMKw2Dngf+JLzFNHgtuvZiv1MglaiXOCQniX/IMC070Bw4jDN
CWmhht0ljQDGdfX5uIclCDg3An9AkHbby0jlCwfmwqX1QcPca6U7wWghvErrnhZoRNvFO4a69GQZ
EEeEnM55paegofcbUUgIDOHWWDhA2s3NGyzo7Iz2hgelTEIXIzquyrls1AV+SxqWqtZuuRQbxtAP
19lRvTIL7mgIRkbXJzsPZcNzYl9CohHaXsSqZNz5ztf52RkfYIQdtmPRlcp1NxUuvwPiIF0c+q1f
JjbP14bF4dkEmrW/Q9liBuN92pvJhQpUCj6kEUg3iDbgnJ5459/QW5F4uh3+MYAMQu9PHlDkDOvx
YpNHApD0qwO3KEdsdBOShhjbVBA2OZmANkKkleiuQqXyF+9hWQpG1i+zPibhXVN7KZBu/kHfXJ1A
ejVmW+5Qs5Kou/dny8ZQZU0N6cu72K2JDqPJW3ju/SSpaotXZFQNyJuZsq0tLiWjOrSDh5uuxpn6
yRIFSMGfj7HJgfilH0ZJvQB93Xp/ROIXorU+hVrk0lWlxQnDQeKVSrZZLM4PgzjldhuYjItUILhV
qIWlL6IpbqRdYT/SIoBDzRmEUMIqV9mz1rRNuXuzo2Bg9Qxj6X7/efpzoMWpr8smUg2tU2qDoP98
bg25GgneyIiKX81BjKel6o9yj3LNmGDDq7ClyCmtPC5ksTUjRIfLcgV18E/8EydwRs/vhDkG580J
DtJmXuDHgeshy+63bLlc7GsSVUJJhjwANxTQ2+4Qgjx8n4oylvutxg+e+tDQWu1JJVHyW6O49iGQ
tdRCd1VMrtoKlzFEkAuGcwW+XfImRRqwFlZpb6QewQx62ZYnNkWdmd3Ua6Sj2hyUUOltZS0HNkUb
c2KzRUyuwBrJq3crEwDJTpQTgFse9v2WULMfyj8OO14ytkxBy/7ad9EKaWkvQSENyj4gXVotoaee
btb64U6PCirL0mGbka+tqZEtXmtcJTPWftSQ/KKPTVlkRPBD3fNtBl7oCLyFiyJW2oeS7a1X8fmc
tqvHW+2eUjHE1+wYholu9u2VxdStfJsIr10B5hbCgH4bGYx6ijGh2NST5wFq7gSmCC7SSIrrO2at
y8Zh+1Rlf5Bx3YIaLIEDCr9il4UvjrudNHaZv+FCXIazF5BtBJSTAQELK01PGJlvqhszXrnnx/l5
9NrhLD2PWqzhxqwavuJtgrNtC0etW0cht1EJTYf324ukIaIt0rIdMYdiWp/mSRxEyjnFeBgU1M3D
CTcdq10THz0atMngPNroYj34mfEpqW1bq/whFF/LJ4+ZckTDe/Ik9TMj1/4o37pWTsRCAH6npQ43
meOqfp1zcYuIwxTDt2EPh1mXvxSmiSpCTPfsXi0BQTRPF7b6J2n20IcIW3ophKYUp2zcMzYwGvY4
94W6kt9aq+qPDBd8WyZCjxMDrarnMimU2+yArceaxX5k9x/hwotnKFLPpUHtB7a7EfX6LYV2Hjtu
gNdJbUZZuB6UD3mA4jLo80dRL1VUjgpBN9wFyI4YkBHyoimUv5iTCd/tsILkFjxPE3yb6z7va2GF
aOyAQNLfKv7A4N4AG0Qj37g5A9UvLHxAKxt5BBG9GA66vxqxPWfBVO+L7pXLXufh97lRRk55QOYD
HLf8y8Kl3fMj3wGmlMrMbTCVk2pp1pdaaxsxcKTcgBB+NmCRW5BtpxbZ3fpeqU07cIU1COaQoFVe
s5vDLmFmbBeAAclrcDM1cD0dAVE+yfS8298hb9cKu5YaDVNicV/iSo28ZzxtNWbgReeGCaYgv3y7
dPlbqr+kSh4LDudO7OLQYRblwrPvExwwAKmEutnD8aGau7maK8kILqe4jV+j/HZaa1BpMayLHBOs
jskTgnZptvaMLyAXuV/GQ/UG0FOsCgatixoSEM24UbihOufaQNMnv69tTqqpa/ifBPeIAjdolx8t
hJo3Z2/Bxgv5IoFBpMwByPK6gz0PsuWPkirfv1TXIwtzgUaPuj3fO8NmnZv2DNHZl3fnPlGcUD/4
B180NRFjou6UZPgmPLG+q9EuokbG0EbSxurwQjpztvdL8dgmrsu5WJRjVdQVHI3CjWG6T1GI9V0O
8tWuJlDScto5hRQNZD7YAgSBuF43MfAT0aMWIgsB2BArEWiX7PN4fqvgiJm5Xg/qyagdoaapFYHD
lIib8dB0zkji8iEQOf68KxBKge0aygfERIw0DaxXXXlkUjQrWTifaLYupOIMwRHtFHXpu5SaLuDI
mcn0noME11svsbPEcs0bCgLtC18jdMvu8/mIyNidqjLBA1YjjsYMWqV/c9ilqBHwv96/TPLhHqYA
fj+QPfzafnoqaDbmYUO9D+fhA7aWqQdODqIoNysQbP++mj78B9I4z5gjIQB8YBeFNc4dCTwq0R4Y
uGitU7KPXw0TRtyKk9fOUj1soq0GH53BnfnadXvX27hm9m1U4252x7SQ2E/M6dKfOzgM4gk76Id9
3hL9Xtea73AumTKfs67qIw22GY/3CFtctRDsXsY6QeQhDhtcYt2feRTPRBf66MnTDOI2xSmV8Kts
ZO4TiYC9Ne/qH5M2AUDO6KM0vBkAFO8OGwE6/5DQeMRCzc+lnef4CcSAPX1aQhUGL5S/0iOJ3dvP
7Dco0oGuCPM90AMgxtRt5QIy0z2bihcx2URoJDI5YGhNBiQ5lBmHp56VhNJ+DtUAkjoK3FCIdiyG
Z+2b09nzWvMtCIp+zD/FY9T6QTRvmGy+RQgP/jDDxS3/JcHGagtOmByWBoRAN+gZR8EtjBgCda/y
JcWbQEvci28f0B98gKKfALm05Fs63KoI4rg6vT4l4lEnGLtf0xtI1+R5f8VuFVb3utuCkW3Kckdm
EG7cuKK7hmAAu/bEveReugOyAR9JLu8T8jdXwTb/Z4JZWHZRq+lgcl1Y11+UpiMaqnLQiA1GOAFt
S5UOdY6Yhh+qbUx1IMX5mVpQLXCdWZzwIQhJDQKX0Ve9CYk9Sia/dltI3XxiKi9rY49kzc6H+lTN
xPPVR/c340MS1Iej/mmPvfFvfaTNAtYe44e9Ag08cmYOcUbja1VYCtg1N2AQ0JOXIdA2j0Em01t9
fnDZ/NglNjDmGdlOmv5A45cYJEZs7LQ1itDnb83owd3JQlIOx9zQiWhfe8eWbTmZ/WqYpzzrTmRy
vXj9/atROzC47vW7RLDtyf6u3QFJZO/6zSntAEDrYTdfenxQqrQFrDe2CCIrgvrUusiYnYm1gnkR
hCIYH7K87Hx5AMuLIv0F7bHnO5uqYLAT0UzgnOsAKEHSu2HF544RCiDZ+LFa8+JgOYU+umrzqUG/
u29v/KZ04pGL5G85VKx1uHP5eVL7/BOZd6jXIVF1e5T2MBZYv64uG39XIL6WGHfutFbNtg3F+C03
1Uc+gGnDo/PdXouJYArcAO57+m2FpP1ejcpaiaHa4OriXF801K/XEZv0luF5w6GgJec4qy2mKXqW
CRgBaeONiczSpgB0JaAlpzQjY8OO4P7+Mw2+mMojQL1uM67NA9PwrE3z1DLeD4CskD4lSdrfu6EX
kdVniO6UmPlzDj/aAX4i9Znt4wnA391hg2k4yfejLK54wvlWIqYyPkO+v/A+Kch0O67PsXP6JcUs
Z1LcZGFFQc7EqiYxunJX2agvXuAZzD+wmHsdguF8jzxXALAgnOBrIW1jFDETsZOMQP8NF+rffPhK
gsCrI+eAw1HzvHCiNC+/JuHcP74HOc1+Ab8GYVMCE2nuLoFgMCZWgXLH9Bxrl+SbV423Vcb65ZP0
Ofu4kSGrsYV0lDgGiPMi4td6Kmi/4FZkkG96XhNO5+tMu7d4KCEtgSb8pBjgDChx7oQLFB4ffUky
0YxfBfhuS7MvNM22ZR84faznuaZ2GDeL0a6FZytvTqgj3FmjBlMze+pfvviWLcUgITSz/Jyvw6ec
HUrMllQLpSw8d3sAV/SHAwcBZs5e9DdcxvuYK6aJwRt+/sOgn5D5TksQSVMKRly6cyw+HBnNh/WP
nOpkyLYzTlJc8ejrD91LFK6K2ezCXlrE0pDzeB4BBUrSVnnmpqP8l/g8OOVshKuurx8rvIdqc+Lp
k3F+XkyaWKlDTZD0Q6FaO5+sYriiOtRxvEf7Tbl+P75+BGMrZZMEu39bLNfQdGLEmEq52vM3hV7C
uscFnvLTk1imz8LOC4KuCDrizqS2Zq4UmyieB7FIUtBYCAdCvfGS2oUIBoATc2SayyaaiqlHgn4w
ovWLnTRiXhbh1D7TthhT6W96HAqyr0qd0WZh9vW5x7pBxLb09y6q+0oINm6ezALUcqdBYyiHrh92
aWKGctb2S/p85PVN5ygbSkwex1+pMtBKESg50KNFu8aZPnaANV0m9KLciUk2GDZo5zdZkNV6BmlC
He3XRnqPrYogY8pH+JVcjbm6MEzX46myUBdwWW0lrZ5jRlZFEOMhJDWMmMJsi3fNeDJxvmEso+ed
bX1RHHVJHd5X7BqRBRi5CGz9I6lj0SfN8Hd0VayIn6o9rYAfkBMmoFDHnngslzIAegq17FDFNAQ8
1GgI7FYfuKV4xlLRXMxEgYHFkmqs6QVqPKfAovB70VYLjpYJ8jTdyxz4MXIFtyMLB+VBqh9dpNEP
5/rxmZRmv3mlwX2WuY41e9nZa5kbPcxu6hHoVLmMPL3IPZ8laiBOrlGruQ2SKz7rfA2gGj+vp3Ga
dKTspYyZY2thlKctnNWv9g7083WRBDW4BuKlLX/66ESB992864HReE3w8Xksls1K6zMUuPE5bbP9
5lKBxc57L18Qs/jBswNfGeyVbAgK2Zr9NARSVi2XycDu0k5kcTbq8X8OSKFSq2UixNTJQYnvqmdq
egg2DJujYjJ6kOeNXxLJkSrQeRMjkOw+dOfupmmkUS0XXUEEui1rSr5JCoVDCyGkwlmhzUMEhkqA
igRKF3f8g5SRRKnX3MtvQvQB1DKk8VYVeIqUG2o00v0439AnI35l8Eya15FlJ4CKAALXkYufAUrS
/A6ope08UvYDjeJghwGW4DWTq5AQWTlmrGV33rLUpP2tiPLVdoG7FU/b/oqV7ohxxLcrbHloOLum
z6SDMls3lGxkslSpf0GU4mG+KhBuOnm9QqyOFGJ2U4TiovG/VjXufsBSRCcX4Ase9lbdHwXVxA5x
Mn6vhWJFe6SFh1UhxZ1qjwY9Lt2xCk/gOXOVeQkP3x6a2UJOawdcize6U2tGcQUXpEGzEoOtfLQa
sII19EVaztmg2bWxQB6vFoDfuWwJiq8wn7MTApG6nEeXdWLxT7fDoKZPlBGKli218tVmxNG408zw
zD+KyIpqGryFQGagaqqg8KdUMepvTk3VoDmzYFMaAAGz2MS5sN/ty7tuibqwOTz9AqAWu8Tez+p5
Fgsei5SPy1WTi9mptuRgsTtCaYA5Se0B1vbLiRMJNTA3avjy5xky7l6aMpfDgO+wP0MXNGhVD8hP
L1esnfcestkptHnRCxplLpnaN25YSsISo15d/ytyHWDf0PfQ0Ig7i7eqwCfB70x+Pm/3Oin+htJ1
i7PtRnw6M5A6BE9M5FOjaDDYULPWpy/tfj/escOOSI0nFERiDiOph9Y3ur5erxeyFrxEs/606hoJ
R1Hsn92+xIiwdW4B1xeAKyytal2zVGV9KdxjYaSTdykmyV0BX94cfUxiMaSR5IGnWFPHLaP6prMa
U/nfMceB8lq+tnvF1pHnEFGA45Cw/3izIvKB9uNikwsKAejDsTWQ4kHvJ1jdlxXG/Xvdvunf3UvR
+slQNZclEv43LnQlhPA9oZc5MH7gss3gY/gL2MjB/Ql0MpjA5CYPkD0KDZ9zVKbM4SOfmhE2zlwg
Qu/ftcOmdwLQz34RCP1ubYYOldd/P5GV0ePHXJZOHKMqNKemiWILEaHz3ZY2IIa6mCEu/T/F95CX
mLKoP1qeDr/1T1rjOIBF6IDJaajSVt64z+8wfAVk6NaZSklkYEa3JKzy1YflXeQH4Wt+SB1R0iRn
zd57tBuyAXQaPFV2PjeF+vbKSImkpwgGimHDmzpOm75NGpSSbND4rgYDyXYdHrk9w0TewWQCq+9q
uORYAZUFrwrUQF2GQ4p3wyp9z/2FIpTHDEGkEC656sLyKAoI7wQ2XGx6DshCfeDw4ysB/na/3VjN
LI4KK4V5PD3p+BMKTkHZpJgRORU4Fs8Mk37RLEVmdvPSkl1zb0zj2sndGw81uX3ZOZC66R4lwVy5
wdORC3dtxTtv+KWVXP3Kx5AesqCMgRq9RhK5XkskPhdzXbuQOFe6x+ypNWf/5I1J5LZFvPzvIpA/
UcBwhDMfp8oxcTGoV/7K+b+wQrby9juQDnopkLo7oAIKlMzketh8IFrjMSwyB8Jt8INAECLfPpav
fVnXfMzrdY2XG1cWUsQqmzMgP90IZDRIF/C5tlalrI90gJrVmwD891pUWL6RJiR/NkLej5mu5l1t
NWGjATUKmAfN8L6InKodFs3suUUcXp4qZyVkUUMVHorcrawO/Ov9ThH2aa8DpqpmjHXUx0Ab1Neg
QNhAAxI6aEnACsok2WMIeoJyqHq37qAiuOFV22ZxE7QFTvn/jI58zPI1BtmWDtYCTaMk+kcYDWrt
9ypbEsGgRxTGWZgopOrtEASy0YmVhS9YYg2DYhTuT5tr9cYYhiGZok2IaSS+YRk3Qpo+q2/nD1px
gzo+UTz2SL1DhS4NVWHyACU1YkW9ixIdIyquWVmd6yVWDnm0BlIs4nHXqYlpMfdugOvGK8K7XCqu
6r5Rl7e/oNkIZjk444G44aIQOzPctOLMypWGruC1FHNitXyD8Wqbi7ffSHhT7/8JjDyf4pGzTH7c
AVXI6UK8B6DNb2T+SJBDvhUCswmxdDZHE9nqDZmw161jRMdkrG4a/LIqauHUYq/+hzpzhBFYxYG6
VHXdvOY9Ir2Qr6nWoG21EzlzYTD+uzulPOpI1Rd+XFXDtelApfdl6lTG5Wv+r0ZuWSgkR6Qv3l5/
8fINLGpuCAFZUWdXxAIX8zvuQBs4Ih6xOn3QsAsz6rLYv9ookQAnrHqklYrwl1szOYMPOtU44Kn/
Z+ShEwNFGaDTMXjpeuyVzCJDkcjRJRzoHWAGvV6w3nCnHHlsRgaCMEkcdzAdLlDc7acNO7nYKOLG
uity+QrF/VCM8C2sdP16JFnr1dJSoQL1PhozZtjeFiN9eaGkbQv4zMsoQegl1bNCOSBcMNN7TL9v
RXOnNK/BtV13seyYOTamxiEa/VSXu24oa4WZEaSK3o0YKPQ1j4F650hthrPaxpjrEnEqo+er7mGX
Wn4tAxuIYLoAHSgn5jikwX2OT2hWxQJhBhAGM6AYJqD3sMKBjYuhvmbkTNSUcu7qhBFKjd+/jXbj
WayQRHrEXYkJSN/46VQ+EEWbp0HtZL01u+Hv/dRMMK4TelXI2QS4iXUwDJKZWloagl9gpLk7uJEb
gF41A+1+mG/W/K1VQepS3xlmuo6TPH8GaN82k0Yjb+FVMfT3Co8LKPf8OrhfZTt8RCzG7WE9bpkN
j719BX4WJ8TUPw7qG4s3LkA05maTEi9Uy30VjquVvCtL4zNscRMeiYaq6TtA2qf/cZT2yDRo2MSO
Hil8jcsul1b4lKB1k1vOYZhRbyQa2zVYdjekD6gT0qrCHWUgHi3GRTN+cujccGxDoVnqQ6UEAbb3
mppj4hxW299FG2v7+bk0sjDCsjcqNCRXKjI1OpxFI24t7EWBiEp9a0IkzLFquwL19D6jB2S+3voa
dwmT8ux70ovbKXGtiKb2Rt80Z1uZBG4NzL1dGYgCCVlVewaJNtouIjTsYmeL5tvVkp/ZxDn34/Xj
6+b5sBKxvii3ZQMlqatA/FPzk0GLgNtbMxH4rx9vDM7B7v84iSbouZwvlH9Xj67f8zdEY+TzD0r6
eDGODsTgPTud2Alh94ihDrLuLGqRH5zXbXhPBOE7puilOJuaPqtqJMZz9CFQp2edeih2WlKdHHQg
YLlISHNmoH+wW5EiS/YaQiNpRq0LyDnIJZE5AcQXLum1IqHIJTPD+8dYdyUjqeCXUSvv6k0z5gMy
5xu4Wx169TWRXuCjdis0N+7KmQXB/XQvfsGw5J7IqIICTIJcwPS2I6yViMLer5Tk0QVvwbbio7dY
G0jrtUxQAZNwWavCg5qpgA7PkAy8oA42jjnpCnNz1uNa8JfvkzfA0ECWABM3/N2zUCHKeSQqNIga
eM9tsZZl3BCz6rwXYdQp0Zs4eD8BShrbXuKSS/hjkeoDSg1KkYXaog9SDwSZDzrId+X1hBeE5SND
PMVXiQo34+T22Sew1Z8fkzd+UJc4zrq0r2g8J4sNcP6D+snwAViCz/SmJmzuZ4XomU+GwNkul4m1
JQdLGNWgywYMCCPLKoMHrsr33ap4MfqEPTy7lHgS+YXL42RTZOw1kUkA1w2fQSjobqvEHWbgjYLu
qOMDpzwvSKxt2sqOKtaKdjTonTGOrD9izLv+WZuC5YAtusDZM4ynn7IGIo/SaVlGXs3xjCcLTMjp
g0IQoGh9PtRohLmlwdZGAirbDMt6DZ0xSFb7XfZ3uA2cX7cNdRJL1yAB+kmVtzEEHHZzFdm41E3g
dDFYr5SsLZEXDhB+DYuQ4pA9XhjgWfx0PSkn4g+NEK2Yz900LwKGxJx3qafq79Q7KYfvKRmH0ptp
xWtqTlctBqtTUTitV0PCmt39whNLm9+eDTjlwCx8hVKvKdR/ai3JAGmUxmDOjBh3wTBXWBy1pLXP
cGq46JKCBzcwoxlYwe1VcDqF6b2kN94GCCoG2KmK5vS+EAAfaF5GsX33ogzFqNxHTHZVsGTXKWSx
DelRH0hBM4Vcvo9Ya1ciRzXcZMQTktZmkt9AmicEKdoVmjWceE1GYaD61iLJZxCRjrRqpl3J6UKO
Mvs5lrCQzVbErB1J/ACCGdRo+sRIyxVxpfYrnJSP85ySv1s8gU5m9bJwX/NvjYyT1werNDl0WAzp
IxEGy9WmItQUgkon9gcC0flLTHKpJhgiFvUZaLT4LsreIsHRYd9X75SfjFn5OI0bqhfdU8B7qxtD
qrr89xIvjUAPTJqi7BErDFpUY0qNXJyPIoLhYfqolsrX+iU0QeUfpjnil/F/Ek0h15tyfu5AnPdK
GuF4E4h81UXVW3gRcKVhXNgLJI6bkGt/4+KI2/ZDenDizm/U9emJbkbf6jQH7bI73uQbxtPpC6sq
T7WTJxSoN38dZF++IbtCTnB4Lkt01kD8uIuvMhl+hYdD/+h88QvaQeRhSCFSK43ER7H/3BQQ9fZM
IdclGd7AVHYBJIcZNMlgffGvs6MAZpFpvX5DQT5QI/7UjwPEw9XFY1iPb7JoyedO2OhLBmD4vONZ
7g06hR1qnSlJQ460DoYMnTSFYiBONP4IV0IyAnJbTCSNVuCe8Nb27axomd5/ArGpaarYX2DOS2+H
0xrkuUj0hHWLg19954YwzxP4Cf942uoztKftHOtfDT7Bgd7EnpuCv+HutQ2eV4a+KWEp17DBLwMO
kNv4qEKHYWC5Kpzf5d1ssBIqxqdDAZfTuyRTlTMJ479lM/HMSXuMnpBqK5/3xGNEB0R6j1YWS/QY
KYJp7Gi10c2tpmK5UgPKgrTJazqZtoWXudL7dX2oPo5fb5roMJE41Z3TzmJZLmPKMzfZb+9ZQscc
rsNyd3+jmqJHitlPp/pDEnAn1LWtcioNPCrd1QIwPUU/IXf6WSdky5LM2RnH6EPv+7tkDOU6nIB0
PL7QdsYmQXlb78nMtQgVBnw3WHnnRQgtXa00rX7XoE9iG356mVPxV+G2QzWQpz/QNM8dFH0AG2qD
9v6ec3rQlUeR4lg4H0iDTlF0aiv6yVEXV2rymrcz/2hB3yg5cgcATaMhhv0m0MeeHS5BWucRGgNB
3uC2hq/K5rA/kpHbyLSDSp/tpsRRo+40BYWEzpZ9PpB9wkl6E1M8Br4hNL/r0EBBJwQwH4X1Ca+r
IP2wRUmwTPmiCRrqXVDNCQNXeIJqzxDmoyjDPKWZOmF8BJFTlnsmHcyQKxusibgsv8SlQxSZL7Z7
qLJMZjKBhiI+weP1QfeTdKfXjhNWZ6yWkOypdcIRjx/twb4r28nYQxOr5OKHH7fEwoxXeMyUnWT1
FG6Hfydgc22v1vg/2QVcMZ7zVNG1zAdKGccM3t94/YKRiE50dlD3etOI+gWOJlpjDqxpeIBjIuqO
OcodFw/2lt5afXdPMnVNDgdv6c45Q6HNKymovTsRc2tx+JAmigPI4eUUM25MKlCJ0Przj+lf5fbs
Zu9e3vfbdj3YQKAXR4jl0faN/eRcD1LjDzH1Rw88KluzUCwKJwcSP67S/q6kzKhmvzy1NNllVMLv
c/S/NAdwN9bH7QUd+18NMnIDyE/AT19f1tH3hbeXf5tshEaV8NTEzgMM5c2Aqe0+r7pCp2HCt40v
EnQSPlrZiOC2T7aHoL4ajGgTpGZRYXUGLmWrXMcFphly2QXRi9O1yWSDMOC62Qtg9WQlB3rSUgB/
G+TvrDphDav6coXfy6ebmDQ0iDEAkhTMzmY9g7O9iyLXXUGbRwGd3gn59jdhhwIZi7y4wInBuKwl
+YniUFvrQkQM6s/v2XGiMuSRnnbiGmLO4h71dv8ptK9Pi9CDLM5YMAiSB5kUBHhHOzI0dNWJge81
HJABi27oSd0sWoswxkkkQJFLMBnMpbmCdneAEb4St0Jh4HCwd/kQuLDaUAFrovTVtaq8wQaSZFe1
bZMxGOVJyAcaVlEwWRGTH4IRX24HlgHo0BczdvAGDYbopQPC7I/baiOgUHbkAZ2tLGK3Us7teV8O
cz/d8BSviMX5T7rtkxVGpRIOsFrSRYp5h/doTD4P5ZluNiQQMcT7XP9kXJp6V1uQvpQL8ooTEPLH
9mR0yLZeFPV+6L5lKyh5rP1dHbHVwPJFonsa/Qvalx3RpJ46cKRcdMhiJUG80Sw0JL6pY0HQXt7i
yjMsmNhOaMDDHbbi+rGMkHccBMCWja5GKPCAUs1H3O9PzZllbh2kydIDc2UpRHIw4HGqMWPx/6lw
al8O62ls6hk81K8R3rsDtFDX2W/sidTE+Q1BvsRSQmT521WUV14zvXi4tkUKS5L0gUHwaAvT1jd8
kbE0LMiVikOca1ezwBHkhyyn+A5s6GG24au/kfcdu9A4BPiKuP6TRhecSjgyPgYd6P8b2YLhrHQ8
upPownBvNz4lEDaiIPXjTZmhC7yrLina68ylXXBUUbhq4Cp5rp81Vp1WAtw+Sl1d2Jh3bR5jXnJM
3JT4sAgMeR23rASsVurOV0KjBgeJJqrfcxZU3Rf0Nwwoze7AEUZ3kWz4zIwZCBZn9AJqKjoCms90
bkfB53r6awnFW8TBr4yCXUEC/4W+7QiSfsMm8NB2Fr/pD0uQA55KslgHpmLmL6PtZ2s7INMWRtDo
DDdfW1lBxy3bX6Yn7StI9czWbDCk8a39yZ/o/0HYAFmztzQIcmD+J4GN+AD6Bmlbejr5ni0eZJoh
D9x+IGOfKeava1Ko4GOoFLx885jaMLHD0uUUA2ZpLWMPdORNeoC6WoIGM0j78Xy31CAJp3YkB2+S
d7YBPbASjV8SFoAaWUlVvBAKOGSQN/CAvrjE7FGxUsmT5FvYnl9v9PClC3ajmtT5jnz8aNOOQhy1
KOAJXYrsK6pWy65PTKP2N2z0qv1Qh3PImbuECTUQukdqkPDOvzi7WdG2YlqgtVLnHlTQfzd89zZx
Cb5VogN5MtB4e42uclsdVYS9Hw7EF/fu3SITTN5GcMIWxSQZ+R5uhptDbMtCrhmY4uw+QbXJqYD1
7G8y4yeJm2gTpinwyHlvT1P6HR9uTBnA4bytSHoN94Ji6l2qtWop0lYMrf6q+dXwE3Z3jl7rRSCt
IaLcYwx9D4mDMeq1bmNzFDqWSgDO/hymK+L2Uc3/vIGE29FqgBuWCx9sPQr66Ap6sMhyAXd3kdjB
U9xE/DoXDUFKq1Q496FAGP8afqWZkgMSy4YZ/Dhztmi9rn27nTL9eKDsg/wL9KxMbYF1+16BVOKW
tN3h/d74M0tqg7G681E9vGqJ5eNv24nWfMJjbzorOGiG3aNF+KAhRNqLLMSZF2l5EemIVZ6v5tTo
JMacWLOgDlYZddpvpDqRgnKtALtD0ayoNb6ZYAsEEXN332PoQaX3wON0SEyiucORu241wGYYS/Oi
98qpIBGICw+iNZj6uB6tVDwOytgdN9Oc1DUlLUzpP+1EDQzn5P+zgwn31QiuWULK8jucReQobe1A
R0Eq5DEJGTd3ktI2stlZLSAyeX/vCxMfK+fb76G1+ngipt7Fqf49ZYhy3wMFbVcN5Gol3Ssg2UFc
wlw6hVtSkkNoshy6Xt1hYzK5VNgybTgA4/x+8BXAzx6BL1KflJeH7jOzWS7YulD50ZztNwezRThf
wYMx5AqNSVTD6AG0PMrSqLjxPQCmS3UxQ7hUM37EcXPmHwoelwj0v9lyCjCoLRzySSq/00CJDiod
kIWpH2b4Rcv7ro1+pJoBzJ3HOLYZjU2S3sI1DGCBJOwFxMu0LszPBbBBSiB5NUcBkjrbfFDn7zYW
qs77EgLW/zILzm9y752/e/FMDukvhfoVCSuD5vKoJdanq7lwrR+SvqQcW2kFSdMPkRJK+xyyu3pS
VgjmS+Ari8xzHdy9tAPCZ2giu8Vg3WpshtjUoyyFzig8lBDaNoe7SzwnVcBCfrJWx87d9bNPQ0jv
nJX9AV5Vpg7v/66LWDmEJL3ce/EFGepq1RYBv7DtGCJZt33jFAF/vORr5u86jjJL2MqJKEK6AVdh
TJZYb44XgbIq2DHZyMSdl8mJUq/P2x3LJe4v0uTt7pA2M8d5+QhmKxLWejZIL4d6YnQgTD6tLn6M
2Jr722r+9bEHbGKnf61JRT42Mb2SR8ez00JhDzBVx/Dwrkzanri8Tpjr98ZMdPzVmdBvBng4Iw1H
2oVvAwpQ21VCF5KMYCElhRwUH7NzNbf211x10e7MXA8+tgqzlWS4s8lFSyCfj92DcppguYMDu77D
wvlpFkWKB0GQod6q606HTxmp8cvkRP5z/QHvk7BSEK9dxqT5PIfsRgqG2PYToKzGF+DU6WTdIl5E
vVP/2rlQBN0i6pikuIbhBLAqBGaxqDUoPDv8L90fMdOOv8Qlt6r+Y68g8bp04EX+N86o3KWHeblF
EQKwnaMZQ/GQWPzstWV2HQEuQw6ERCKYygy/C0Ra32oE2dTiUOVMMbc0slwPm4ICT+IMpxYt5l2S
kDaI0WOFYYCWFovqO0P6+3py2DeAN1LcNHQPwo+O8IFa8v7nnveH2rcFa71zhgXH+jtVaSC5dBtJ
NCQVwfh48ziZha1NBCIhXp/R9Kadsm4f/IqkkLlAgNPawcxzBAT4vEcgZPRI5tb9JEZu73Rr7JuJ
RqSv25T/adO9NjvSLeXSclTL379epoTV8w6kiG8s2mzFv2QVO8jxf0Cc7OKZX58ZNrRSsSaxhj4q
2yKc6GHKByuaxuqvi3dEVcs5e1Khgz/5AHkiONZphA9HFRH45kOH9oxFhG65A4QqLLfU6jXNdMqP
Q+DVMVSLSwfeHCPPuw1AM3j9Mcg7yKCCzHEXo1qqdVgaTxb5E//P1zNv19hIRPOMeXN+twOYi2cs
Te6t1ymEzZSl2xmZ5C/7CWvk8iqP18yKhWukmJSYST5U0UJ9xKIghqn2jK4wvAuwpooBox7NpV3U
mocTM28y1ZOc47GXmrPCT/sg6mu35jLdLxUsaPhFpkqfbPPvIJStlUzvoqB0GdsbNZsS7/4CoMTI
R51TuGeYGd2Q1XI6RUE9ycTjwl6xjlSa7F/iunBiYkSkkLOU0SvKs+SPSoE+8UFtbK7dl6nBXM3R
tY88DYjFJuxlBPtdIeS9nM0thXathcCuBxGw/QWWUuuhY+tIw/0zKd3158A9r2WTWz9IhEIf5Qld
vYuyi4KogtYlhzln4HH/rH12Rloo8qTJFSWQsiqgNVTV0aeaQRy6TRZ8XNVIBs3CKh/W9myIeM2p
qlS1IZfot7kJbJ1a/Spu3alRalxVGYZxqOVMkbPO3hE/Ui3ntOeAISAPAelg8P+naS5FA6KE7CpA
snAJeRtweEZN0ddIeGErDYDt7HuQ558kjjLI1551aciemzjyM+SV8BVh8piLKBPMfu+63Vz3IDih
i8oHeHpGh+sRRygaKvCy6Jl4yaAT6deSfpEhbMXe+af9IRyI46sXupUuhcYAdBRSs/Plvg1M6hLX
dE1xT2u/S6T1RhM/xz5H9epGwl+7Jqm3JogVNaZ9lnE9vTXWhFtP0aWvSlXOw/Di/rExQ4GywkwF
d2iP7NWk5el5J9JzpkOV9csmvYOOSEtO7TktOZODFquqxjFuxSmk9S8+WobBAy4fWECfonlIT68A
ieCgfH9auz8WJvCJerkRvsKlMVWoFatNY+atzHbKz3CjcrX2aAm8EhddcWwhCVIHFwZBQaUVesiI
eZzZIEWNNk4G9Q4bY4AQeWb2/Qd2aDDcCHlBgXsr+HFsFWuuRGtgKt8aHHX0HK0kv8lKVv1pi+Rp
EmahmHvHCdOFcTLMcydB8PPqYgxZDhUl4WD2Gzt2Zn1chOG2bl2MFd9yCN6w8uS0qg8ovQPxWxNF
eiSqD7D7PedTS86/MUhK1ar6+WAjxx+yRaAjni53JatKLjV2lETkAcx6gMs8DEQH4tmes1LgLaVq
fXGladTH+1HJaREaR43MqDN/fxlIVbiFnGPGL/I9llHu3U3+Aypn3pbH0CmXJQYEJ7dKvfoj+VMT
wmH8hiuGRg1sseOum44gzLRJOs6ZCDNDbOPJiQXJaQ4pyxJVvf4mwkyOPqL0jO+pe4+WtQc3IiPn
OjmQVJujyJkEEkeYS9NTIDjedd6BgFP4Lrhlc8Rr4dyCTaR/A4d6A+wHZdp01TsZ0O3AaNeI9gqR
gnNmJBMfR940IXT9Dm90ky68JJYydcQRKLOcTEfpAbrXQIXBKEYyRsxDmwgLC0DGpOYYi03EHIsA
v+nr9Dg/g/+ZccbL9f1e9h9wBHcWk9/jZ+fwj6GlcpkSI/+QzGfLukIk9PCSPJXDVskp5O4puYDi
TChpFnCRb3xCzNX7CSlPDckFmt7ufRv2EorltHsW+1q58zx3MteDxbfci1q8/M+g8IgKQpZp1Si1
rL/c7RVkcR+mjViX+SQSpwEugSgqzv9a/yuaV5SN+jB0AUhzAejruOugd3kXw8VKidQO0nKZstUF
RwWVj0Y6vUm0in/aMvrfslMeBKBTLd7ISYa9Hc9sJDQ6OYxtDUf/MjB9l4VyQHsOpqQDp/3Q4U7n
IqJimkKy3TU+P9Z8wEFjkfIacc79M4dQS5jCG7xrdw4P1sjpLEbWWNzUkil8KaHOaoYDg9ruMjtT
qIVKB1M3CqM8+J2cV9ZueSCPk5XP2pPaAEQ97dAqOV6jMvm4Y5TZhx2aJlTzvGyoyZI8e6tobQml
RaHHXOhRgMY1OIYnUXpSMbgpw8O1a47/TV9TgapPLWAbBZ4tqUhKdpEYKWo8toGfdjdbbiyRQAhO
hTNK9g5pZkphl6IYtZXBpOmtzZqYGax3niJ/1g5lfB3VoRHlqkfrMLb2PHcWhUtx/126Qq6Kq0+t
EG+M6t5gXH8CZfLrRDjA8BiYG84P+n3s6c4OpXqXl2zHhj78ARA2vNGeeSpwS3XP/LpZ74atl2JH
mHG0s2b151DIa5vqtJpQ48ib2gvFo8GAq3eUmS8IC0uAVoX2wuait66KPk0JMQs4+suyIQi4jjTb
TGBKIFm6ZIEfwFZltMJ90JzI36MrM0Wb+yxSQ7UzdSJ3uXQL7iQlIfdeH7NtIeEaFOulGSASPcxE
RKASSZ+7zapeQ0HUpff4EM/NzFyssqz/W9lp1dF8CyZrzym8pBVOX58ny6hZ9Y824JLYDkF/6nC9
k7Vw4W6OefafW0CXGFbmNWHz5Y6u4X8nYpZE+ah2UkuXsFqfBT9YdhCvBHq8Yx30PqiwV+/DjQL+
jj0XXH9uk1L9cF1nzVbEoMhd9RCA62Vacr+I8A6ClSnvBsJa3lAub7bY4Qw7NqO1+AlC9S9B6XCQ
GLZV97W7KSX/gChOCBKZWwnNLO+Rlvup7phfez77QHJ0iSKSjz/OOhagc1NzdWhfNS1OtlBYFM2C
R0hye0eO5x9T/1Q0L7jUhwgnfpVu2bs6drQBVQKsRcfSy/Xuv8q2C/HM1jGHGJ9tFKYwggFmakPk
Ekit2FrAan5gsGCyBGa8Pu5APhDfghYsczj6HlG+YBh3bWmn4R0mdSnqNATGFlRFy/yEFI6xVBoZ
8CLKKqZcuIsNh2v11MKVIuOC/TkneFLiQMyMGjQzscBpbXgID2NH1om2zaNeag1FhIsF3YgNwAHG
obmcvVz400k4GaPusYEK1+ml3gWtKKWfU5gAsr0wOY69dU7z8W3mKgONwVRy04TZKWq8TNzEb+zj
mEqXUdbuN/K4R8UHu52Q0Jhorxa/NTFTHFZQ7TLB3ItDnZ1+9yYlQV5iSy5G9DNi3Gbz7K8HaVPP
cEJcknPnh+uELbgqhyQ03T6tLc2HrgaVMm7M9VAhdjrS6nD5QovdcrpBzxYWgHFojEu2ecPwepWA
vBZJOS8i0MRFHPGoyC1YusCp1mjpKZ403yV11zHs2W/u3dCpg+CgGG+DdCKGDYKI/aNWfSoalThI
k72TNH94Zhj9v/42wvnfbAB3t5UHjNIvImyr3tiuSAXEHico9/uoCKwVngOTlKaQTOT4ha1+aJtu
OFuH6bJJsRRu5VDGouwar+Bo2dmsLom7Vp0W+rFU8Cg4FFX+YfB7u97AaBVhR6oPDrPkrrZriV+9
UX1kL0TzRsh86OI2td0PSrvafvy0PQT+8SO/GqM0GZdbLuA8AMUg+TTMP5GIDlAWUoLe5kmIKR7t
Ed3tD2oJjqtn8i1NGBRgp+0murCov5kVK3nO7Spdch4II51FMRvfYA3LiVfVNuP7k0XobtuJMHG3
xXyuYnCdeaIR/om/X2Hpdb0UjC9EU3QvtRFTqRqQmRAT/6jzd87cR67GWXJXp+DkPgq64OU9Hjqx
lYb97e88vtp2S3yALXT9AAIKbep+6mUknaE2yHfjzmaxo1ApMRqMlm8yw3DrEv3V/Dp6wim9BTOE
y7DcTRiAxzvJYdUBRGbQr94C66uGQSaQxbaLtUEdoN52itauPJ17Hqk7wBhMa5XXtzZftdUesJYQ
WUVirY62k+3JuEbQGHiaa1tt6i4CIr2IOt6zJrjQ1XvB5kz/qE/aJdQzJNFaIiBKg52z+v0ciDMb
1zEj4LQ1km5DmgtI9S5mxl9jeJM/R7okZaoqBEQAv/yCNGZxqd//U3pPEbTo4WbC370/yFvzkqZL
aflD29vaKFUuIcJQVc1bmgsQooDPlkKD0bIfqirLKDlfqYAjNa1eP2VctCFSoxkvX/czGgWY+gAF
0A6ZWa0fGWy+qz1LvJUtk6DEbwRzrACWrlNp8mx7/WtJGYnk+EgiHnL3mTNEV0eKz6VeFjuxEUwY
gmDCduXp5kWruOqSq1hfeZdnYmIAo4cxQj4oZRdf08wSeZtrJaL/hRkmvXhSzhU2SDfL+pRYkC/x
ErQ5F5Yk3iWIVg6PctCXdfUNPas8TZ8s2pP75auZO0ZuphRxqTO0n+5b0HA4Tnx+Fpsy8seXj5UO
zLXDWN1OLjoHQaUEr0Yc07CJyxOgU+xT5PYxC+BE66ni7fFFCIKd6VnrmV2bZ39ZyYa93i0K6Elf
lR7zBcWC9SPmKC1AOWQ2AiJUzkzEbLKxQK8SA/nd6H66tso5/Wx0EZMWAiA4snpMIsYOTw4J/QQI
csElRQFdFBvOjhJTtUvskfZF1V9OuFs3BTBIEOXL9Pb2s1OlH5NH1wce8PyNX5lPUjPiKXsJiiAj
l6Fh4BJQ/G2kIwuOlSOmr81CuZo8obi+NzkfvbFa3xUHg83RrTSYnZn6JJ1ApnHVluljy7wSqriu
onFrjUtU26YEW/oKHcuJAOIuxMdg7/K8buMMr67ji2gLPosXdBS8yGS9HTgUiiTLqmlRLZzV45zN
0v7kaWXC23sHpSzre0BBIswhKGTtw4o5iQt5KfwBF6sTz7PuofaukHo/RRcttVqhiSh2ocWunQXw
DdxgfJSQ+Iey4YKBKKFw+C3BjUsFEmBSm+1FSEMfD8xiHpp7xYKEbNHCgkIlvu7m0j+OPkmUhjjx
1xAbfJtqRRnoEizeDc3tKn+hhG6d8mG+GxRgYExRv/OnXlyNewhtKJVe3ZsTrifABBn8t6iAIFtA
tBZclCzz8dBIGmI4RD5QqH+XiLs6B610RrthS4UqAmMmSzZibtAVT7LoyzLfxRurzWuBD5buTCzb
8rANQGd+drMjw1Ss2nrTiKqnLZr9O5ikFqMEIN6+kZwCFYoCdxJ+upkTeROX5VYf8V0L2akA1Cy9
cCmpRNQZgeSKEpJGZA3mBj3uWBeQBe4PgAXWUUdtp9TW1nSPnpv/BEyFSYahNebrA9iI2E6JeBcM
LfZXu+wYKHRhtwcNq+HwwBnU7TcV96n+XQVxcSAa/GYVhx3aObxzPmqDzVUj4VyortpI6xP2pEWA
L+DFS7ml9GxQ1X6fzmn6UCRZdDyNVaZLT1Kx9O/T6pkpeOOkkOKfCT3sV+EOulmA2bgQZyBm1DR8
P56LvJXmJGZB0/mRxQX74FVKbUlJx48vuk5EgnagUbcda/6sQJv4jiSR160aiiIaw2VAONkcfsUI
Nz5DBIjvv4PcG3c2/WjgYxkcKKLwuHRuy34x/qO+l2lePMM20BAFq/FjcdfTI+5ZIjyJQi/cH/WV
HIrwT9+uBfFNhsRWg+EB8v41RGMscMJzvM+8r0xuc+bnFfH5B6rnkkrXywGVlAEwNKjJ0blIGAX2
hxXJaO+neuQ+YdNHo+aqO3zjLD3BaoZMG5lfNfgu5XXZenlkagJQFjfEJ+bCPO7zrqDH8Gyx+NPR
TXS0ggGNQNAg1+e+S600tXylftA4c+8BhfkygAG/HTEUMe0zxIka8m3xiaE0o63dXVNHz0a+xI/d
KisB2vRQg4rDU9WEJEBeyDy5+dPpeX52Y7cBnIzMIWEI5mPM2g6EhKv0U4pwiDoNaL7n/0dmkASt
6mQ3vqngqCdFoIGMdwnUgksyaiYGh9sIiI2YlzOq5yqxOTm9BCtm6dB69dpN6ppeJj8rlpcDeqCh
MJJRoWlQiuWRmO33GYMh/Gt+l4gAr5FoWds+NDNplpA+PTiI773e80pGDWucMKh1vqgY8wYTsr/i
Y4whvjuG9b2AIjfUM9Hxua1Sohw/VYTZeCo7PE33SdrpXalSRz3Yb/Mcg3BdZ+BcXF9+u7KjrUVc
yAEgSlSoNTnRDnjxSm4dHMHxmRWRXzTcfRLBrwX+omQrDM8LFcCfK2ab6z+hJkREQIepTiNITArT
1nuztVchERPCCfInLbTjdY4cy2xB5nTWoRoO0XGWK3XT9i13ol+S1jIiyx1OsYtpS63A199cHOPe
LZywIfIr6NVrzaPfQc3yErFYtKKt43nQla+JavNkpT6r0oIZpuYSOh3CCPvKIKqYY1KmgV76xJMP
QgBUZfytAQiKcYc/LGG0b59GXIMCUpptcKgvGaUUgd8cd9jzzIb1YI5LzUXfMJljcREUBtQZQ2CP
Y+PUCFzjsX7HBL42sH1Jl0vcFUqO0gtQ2JJU4GYYkaSkDaV5RUwStaBqAoArtpYlcmDMynIm3ySV
9ao8W+kmttxH5czrz5kHOCDSVpdpTY+zyaJRh8jebEWuSUybwbgnaC5ZfxtFbQx87nJAveWT86t6
Y+5Agu1QQFqP0uQL+RpT83AypY3R99zZNBhONPmTabFYf/6yU2X6xoHx/GQdBGb60sqO+r2NCFj6
7KzXJD70WfF+jD41Yu/etwe4V7QXfterTg0MCCVEVa3lklFgc5u12R1QEc6JrFCHXZAOu2FvbB5u
GGVe+w7qJVe5DlxOEToP5egbkpnSbgLMMn+XQP6UoSqn3vcbgFyVQX2Fbl1M07QNynTthtpR1etE
bFgmI5CwUdBPATb0W7tl9//aWcbv6JrRCB3TAkUxCvMaK7RxOuMbRz6LZUOQt4NO2VGW+jwI4gwW
AUi1y69qVkT4iYI2Rx438ZwnPxXlgPzWYylYrJerTkHTLqB8PUlklLUVa1rojN29BBuwwuMVnUFb
1a+yqCP+C+Ea7QEHN1pUT0wV4KP42o5FG6aVQ/m1Mp7pFDEfOjtB2RtYFRYdboI9vSHiglCD1ZQi
HqLZvs6AXfLsaOWH8dKgRhz8xuwJ7RHG6+N7A4DYd/oaSOGYhLX/xjJMqv7+oUjptbjj+cBsQ9NL
wLzFdW4qbeJY9KVzgpABo5pDyCOKO/5QZLZZI4xuveRWF5OupAI7x3DoIB8SSTrpYLQMukR1qWTa
AosUqYWym/MH1C/g6UAlGERlcQohLWSZdbi6m/BUSA9UGr1tjfh0+FnNAtsJIEfXBAY666u/rc8a
PQeWGEOuyAKgBeCTMIuMLOT91XstMvaQPpHettndG84fyu21UXzXXtX8OU9uzID19n98vhcpyOBC
G67eCo+k4JXoY9mxlICRSATpEZ4uWGvj8UF1WygtX2fecE3JfifEw0ZY0Wu3e9vHz3ZEzpZfQRjO
DUQkAe+PKEvldtXk1XqsxakAqFeCY1iLsHP4Hi9XQRcA0M5jeBu081RfXbwVPwnL8rMRWkuzYVlk
S2213PdoXQBGg08bEQAk7f2ldt0gs61ofUC5TnC7K53uwzAtZ6ZsOxIb8y6lMg82NE8CHeWMQM+i
R/XQjAY1Aq0d3TpuGJAmu5ibw4s2y0HesbqqqaNiEcuJjTE1JLfUDKX+ceE0vnu1uh8bIc6UxC9T
ITz81oZFhaRbrkzEjlmvFwtpCJGSatrhYrAQ9H4DEnNFqoX/ggYrrOqQRe2ElvjIvComPvEZGN81
t8j1Rv4B1XHl6+4fOlE6aM2B9UprtReqQCjMQlb49EBcqA/4AyisZZk7RM0dRG2MiFdg+WamjgfS
DK/y5OmyX3jWlVq2LBSAUCXSRfC8nmXPtejTmepKo5SkcKnadgE3eCDcXAcXG9Saoz4BNBeWgMi3
I2Qb3LR4sEkQ2+F735DEg4jFPSGaZp/7ZRfNUcnOyabPd7+DBaaQ0ynCv1iVw7r2I2xvnVZ6J1Mt
00N3VQhiDNTP/3TMsiSvV2tTXuAXr/Z6m9X/M6PB/+WhpcT3CYyQauh1R768WozBRhgOLBKpGiwW
ZqW0yAZL3H7p3cPD3p/QebkgQUrsGFkwryLgsqeFdf6q1aRoOxKc0o69JI6bFfM5HEOXj/q+Ik6W
iX7YWfWH4YTIWfKpnQ663VKtjTLZaYQfQ8S5kZw+1Kr7oQ80NY5M+bf+0IgqDxDyKFUD/tBOEBSS
hO4KCL3zyJuqAs7WB2rkYRkh+rJWj9SKY71aDNjYBp65osVL3s/sGkN/h7Ur1Dz5w483FK8aLw7q
iLqkD2iLKyXpP2kvRaXudsacYDH5yjxh3Ve5gd4N415T171eNrQaBuUDUo1if/5Jt6gxXPE73Xc4
oOB81K7CfTvCNMbj5oO/JyzI4II57gD+bOx71e/24eX9DgZ3bbHyV5oPH3u47+Q29d5Thd4x8QjY
I8sZhBXp0N33uIykGPw++2y7iWY+r1RoFo4qf5IHCAutjAn0E+nHFkCPA6SOJ4DZSNK40JjUdIjh
BH6pcKv5WVYZy4UWTItw2uF39kJdoblRrWaP9A6UrxkatPQVxZOSEXLF9s4+QoiolSf5c3yDacMS
Nx9k+ENksmIkB6Lv5jt9La0Mn/dP5suL8rr7qak9aEB04IaFg9RXSCdvzQCbOqgT3GwSPS3RzlUe
SObBuoNhpP19rRQfonZ9rOdKDq1yjhCy86uiMhOXf0U1wYpJRFUlpRbpkxxNQr5PpYDTi2GsTqAz
jN+7sHft2k8CRxUzQQFTrH87lh56E/NP6uCAJze00V0p3b2leh7sbNJgYPxql12cgCFLj3esyDln
Oavbw+jBIzUKVRbbLkJRsGSCxXwTJijOyYOI24cOFL5KAOUKhh5Ws7+NQHRNo94JGwG+WmeJFx7k
lQcnp/fJft2qIUSDi6n5+kntyvTxQCNk6mJrvp4VMCYjCHchPTprlyVvMKL9PESux+u5ltKYeLTV
Fuj3LJ8kaf2EUw/DDMSrGfM3IGKLCtdURHC16Z/rYrTMbQe0k1eIxr0gLjhSp3Ty41AzEB4Hwgkh
sB+PE9GDjDQM41N/768AWJqxicTimU6vlwDPETfQCTbeohPk4+iFtJr3B5MttWthWxrFaA6rtSca
gUOpnxWA3rH7a7Tt3tyfhNDfouCSvOOM4eSPmojtN7uUiLS0dgP448l77tqrMesy0JVnVOCzuGhO
j+O6pI8ixIp2b3Oq3WwKNljsdGV8PVvRhBjbb1m3B/Y+WSfnpL3+SgYfhsKFBHE+6lEIeZ0ELuU8
HEeGa9qO6T3+Rv7vSBIRmQD/Gc3YaqMhLA7e1/9gn/WDvLsF65oD5TVFlMbOa+bM2Lq6Roj1zM7t
PWtWaPIpitM40slLI7+304Ra0JVBrMj6dcY34eaGYLq8+L15nDePJg+b18OfW5ODVeaGCya0lF1H
YLhF8sMQYkzXiTYb6NseOX76d0yBjJ5M8ec8EpWSCyZurgQ2KZMsyNch7fsHLqHBW4vIEt1tlAax
x1gkRVSzIgpjtFavsHnpkAraCLhr6lYu6hi6NEivPRfUuWVUdDRU5OytIRma/qVJ0ArpJ+yL0A6E
JLGs1z+1Xws+7fSM8rcBYOug0jlfpFgrwmryyCAZ50Akn+PNDpH+22HIjtrwTYKfhgp2fQaBr7e0
m+KdaZdKcNeNueIUKV1MYUYVnVcZIH8ETBHyb4dvVx7VYH1gbiBUhvKSkxW2LxY3868H7GGaV+Ps
BNCmlY0Ra8qimwcEj+EETNQZoSXVykkSuFOht/QmOjUwR7dDb9E7dwhzstjht5ubrso7c1OgcVKq
bztyaedLTvJAHv75/MXNV/oQtAR0uftVUcg9pvw05M8daq5o/payEFiBEWIZeBat+NvF3+Lj4ODL
+v5sUP+VecPFpI6VSA4tNPJcwMRoWDQwS59nHVppU/lUaaYqOu97w9JX9/nolugxySxe4TZFCIYb
OVaC3C0QNJzpJUJpMjTgJs1ofn8KkMIODE0xjvvk2oSe1Y80oEs9nJWbYaCf8Dt9XpUhIy/TTuPQ
jLJW6lPlDio0G7hlVhhct4C4hayeGbd7F6JQtoYohffWc82uEKP5euDq05MA38OARO8Wyfv6B4Rg
N69ab1Ogu589OV45PScNqJWc5NIZkYsCWHiLUuIcLXd9gGaRQo8zKNGQCv+sQs+/AkkpXimcQr8O
ONA8UTluDUjZeyX0pc/F8fJE2XusTYuwtd03zwJAv80ZrzZ4ug99QHCI6/DL5BFfME5pS20/PytR
6DyZqzOKww8nPi5TVu5N94PCxHWLx8OSgr0f0ci1oTHFnMkf5aMDdmzCcjFxSXAMHRBbM/tCcuzG
2QFvZj3Xtb4dTkWVqDTxca/eG12EPovvXyqMikg65mCqRIpnhVy8YNPxoGP2ggk4zFrbVxCjLcql
CZUsmi+DOaKdA40q3K151mcn1qk3Z9IO4dAXYtQLhj/xm5KpNX3MudWRArmefI4EosJ4jlGP3zNo
oQIV/Yn8fLo7HMaJWIYdXjeC940pxJggzpiY/bM8g9AAWP/3UKYdiRm3jPWMxtjrNkHhy8uoMNcl
U2O8j3vJWkgqvQfzEw1HOiZRmAuav0Gh8uae9eY+kZsBDz41lPrRIyf6uslzJRIkW+rfNMRtGCPz
MWvmWL7AOS7xMcm8y2K6DP6uGFVD1EKMoPUQ24Kxk/G7SuOLaKyXAsm2WjGSg41A03AoU7ptXCw/
9xUVuxcNuH5NumNiPadAachM1Wbuq2/UKX/6l6orki4oFMVP8IicNfkwE448TLKPoLXk+zuvm1MF
p94F0Nz9OoDn78o9Ra0XdcIGxfTH5t4lypHapghBh53UqiCsbzO9axpcPsC8UGq1HoNYEclP3bnq
ofxTSNWYbnKfluqjxXwRj+pO3XSru3O3Fv42R1jkM2BpQ5PrntATXbP7gx5x3eIgb4WL6NmUMzNT
jf/pfqWETE9ffRh6qFAyBRAMqhoc1PGf6kOK3OTwQhMGW8JO8yaIfGtcRoh2KObK6DVTB6XkRI7Q
6puHImTP/qu1Hc0y0mJnlhMJvv41z/HB/n66DWp/P2n1eIOodIbuYPaxZDVjIprfqilFQGCe4ond
r8LYOOfuMa6jB1NzIUM65qGs6sAUK1a51ulFeDERRG8rfDUQKni/iNSaQ5ItVXDY2rR7fz6qMEA5
5e+G2JIluPAgraJOJJskNRAFCEywW7tamNgayvZ7GVZqRW1XO+JU9Jn0Ca6MwrDN1B55+6ImhOM7
Srtu8Y8IVCz+7+hTfB+rmxYY8JQwpzqcj+/cvt6tCylxQByw8DWhZJUboKZJhw+bumrP/B+QkMYF
enWHhuXqhroSgj+zwqYcFr9RqWjpNEMHY4ZII2H5bCHP7t/zi7edGaiuO+reQc8HpRzDNMjb9s7L
g9ooHEjDIsF9hibzCyjNgkLyj6ImesW4pcs6HZcd4HE1jjakIvAto2gjPYYTxZPk0llAMDUU5i54
C7qw6jGSNtey9j4shGeoVLtbSSSCmDzPgs71qyivSbFlA8TzcRW7rWBArFEg+IxGZpc4zD/rYZxS
ts1o7o6BkI/VRLe7WbLsCMfoNFNh/IuSERM+7wuEGV7Wqv2f5ViZPO0Z6A1ezwypV5eMOv+1MTcz
0dIymvX/FiAO8068HqGtqd3WAHbcT3ZThKKiinLwpOWK3+/pDIF6BgcEKY/CvQlwHJErY9N/b9Zb
9hP1ykFM5cN8lt4m+bpYeZUBIBQghE0NDEpFkh/0Eyq+kusyZOLIiE3OEbX6zf44iRdp6Zduwc4l
N4yFPYw/+olrLMMRiowiBGZ063IqyAbcXwihQrkQbhQ9Ykwl7Ay4Gjnnf6B5AOPsFTF8zFQqNtD/
m+dJP7yuCRhTrvC4fzWDlnx+cp1YwD9uSVyuVuMM3XbkppxwbiCLfVxK+WiBie705k/XLWTpvPFC
62jkbbRR3l+i2Q/xt7FAnKI4gZhj+2jyKrVhVVkrpCyDTqCyXdMsZkDGFa0M/SpUqaRlVB9qwK+8
NIsU0MkX7I3y4if/0hsWb1JRkNv6LJlfXdxIOdrNNayGwXGwomIc7Kk8xu2IdO4bT1tn9RYlpMhK
Vwe0H+YKBDqzyRFvs8b7FTr6t3oKYvmA4fdbS8c1xASPdqdiswrumKq4+ip+BnpiOTlBOUd54EUA
Jjvh3nJEL3WV3TE7i89iuaLz4uwUMks0CLp1pYUn7k5fkREkEC7P4hB9QfSZuc0CxraoAk0ZD+/D
03vTthN7R0PCPb8zAALy/7J+xEVPZJrLedTRcZP+fYNHbpBHJqfwSOer3D5yiI9jMQy8wnF16kkp
qXYYRgxxZhilkO+QNQfX/cwU9IvI8AXsjcoZCRq1br003AmSc3Mwvua3UQCPJzfmUQCT0OlvM7MF
yVdNpfgeLTkiSHHw00m4k8VbLUdH4ITWWGUzFkJ4xos87DLsHW2SrLTUyAGeDOwWUG0V1qIAmKtk
5c22ALLF/ggdW9F+PhIZ5UJv+cJRq/CYGV6Jz0tDHIhpGIzbo8FNA23lofcPJRvmPYmzpFoJ7z/c
qQgitICU/2t4VqSlovktdyxNrsYCQO0RrfULrCOUFOY2EYEVKDisbm3hEY2Y8wG5STVSL65SkoBD
CP5R4vFHWprOsYDhhxAZ6RxpZwGQXDLD7JT9LKz6SHi2C5UARS6w0nlzVMOItin25sw14vzgvSgm
TvnEtLDX1CRwgrCquiHAIHqZXh3EduuLD3y3hfYhbF62yDhNGDCFHRarjugDESXm+QFJKmY7VJrp
v9Fu31X4FWTyksyfjz2WvT5W8X6YAntTfLy/S+4RTteMhdKBQ7iBjR1ZU8I3GG72lHUnjyf0elXi
Yi4FaAMZEibgna+6A3eknYUqC80FSlvTzqg7Os/DWEERbnzKLwQ5zXogORRuXvvRTlJeVQcloiWV
m9EcjTJ4HHNZnd2IC32eQOxDdn8KLmL5vbR+P9c6ts7hmDTLfsUDOtr5A/Vjag9SZrukas/LBMcK
1fHfBt4D5Kf32EK1b6jrTlLQyqFs+NT0n0ftPHaOUJbaMj86DNpN2YD1y7xH8xYHBUYV7QFjSwUj
VbokzCOotmfEIy0rq07yDeTfru0hnDID7OQJVutIl7rQhYrZCAmVHhHjJYHMlNRHpO/kua1ZciVK
AR+7XbnKvAem3ldrGjD9DGhv8EyDWTqtapUC4aWlOVYpp+3M9MdvSIQJM+Jpbb7S+ymFX/4BDMoR
nMmk1FgCJHJslXOIioyN+I8whKyPHFi/5bxv1+dqH/QOAaqkC/4m1gLcd+tF9pW8czeOy9ITx/JX
DLROzEUvYLgAdR8IBGCZKuuUQ+yTP0KI9aZemlNUy+zxU74/5OPHzLt2uxg51aJS9Gzv0YpTlPmb
fv4+rfa/DyI1+o4MD3+gWV/gPXIXqsfoOAS7jkpnrQkfpnrNt0utN+/Dcs66Nl/Xkekpl8qKXK6o
wLlZY1BOgGN0F/Sw3MWL+7NYkoFTdP8aRZj49Op5dYVh3knn7gOlXw5TVtvTdatJ0uYuWtlDZ6Rm
lobgS37xaYhLNaLsIV11vQLbW4FOU/zodsxOinu6bd6CpHuIIOzQNrPu8cyHUHXJ4jhh5x81Bnib
HIZuDXqNbD51pNnFvtPmfI2+Lho4Ln/pCBM8+RIjpN2obLEXOgIwdNfy1Un+Mn0/LGQrTKEJ3Rb5
9vBATrc9XeDEAXZZsWsaA8XrVPf4GAhX4Q0A4GH8dALSMnvEpakRf4KruEe5WxFWvSWU0dezipRr
yGkIIpfqsUNz1efZf420arcaBPUdYOQYThhbyyteGA6vO3TtksDkFlQoRV6OX1VQHnvJRtdUQFzv
q3TxEOkQKvJrlnL2Jt8/lclW2302faVdLQuHCTn+mNLp8rqGEs3+4vInWv82C9bxnjYj7NJdakpT
5RLMdZ9WWIumExtmvP/lfueig25+JTHfNgGpjH6B7n3PUwlFyO3jAAP7x8BwGSdr0SxR9KjGqLod
c77EUsG2sPOj/2+EFmMjrlO+52vj2jLHr1WR7fYuprs0Z89Q5ZEOGb8MnpXVByqj56MqSB+eqKaN
64v+YWd8MqOoh7V2jlFsHF9mfwWpi2G/0NXLInGOP/2AQK9HXv2JV3E3lAOd4ymCubuQTm0yDxEj
SA8sS3y/P8ZsrNZWFrF1gZHDXRI851rkuU0UI2dNot8PYhjzWmIvC5bjHxZhcpigaoqFO24ufhDY
/yjGZKN9mtTDs1knfvaBfZP2Y4LZaBNhna4izqBLYGXD9KYk5X9I1em30P7sA+LMgDtdMVOwtaS3
VZ/rxsJWhojQ2l6n3lchBhRmFzOT5NL7A8Px2NJEqPt9fJt9aeocGLhNLzfVrjB69QatzsXIeZz/
sP8zT3dpctHLWX7LpDAQlV3hX6RzOk8Bly5q/KIHEtuAWVInxEiNoJhU4eg5vPxMfhyEzEJIF0ha
uVrpdh3jtKLExn1/cagWyPC4PEiOEx0YekSSIs7lccDG3l9WJGbLZdJjCJmbqDihrlTmAEyqEW4U
5MvTaTdaZim9Sm2S8uWpdJsVGZzMgrHCOyDdAaEdYivzhOA5ItQ3PcZq19VGhXJKjicwk6gZDHIO
sA4UKcIpPwDR3g1sHixKTdYMgglI2opB0xGmarsRxYmh3bgWG6NwS5dzKIfIRUOs13YNIFfetBrG
PvovwglfdmZnhlO68jEHIJPREP/efB6X4t2aSKLZlTuSt4pukT9kABT2p398Lwz+vp6NRDKpGIvR
OEq9WphPlSAXqc4BNQymjuKPbFUb/ZEMCklTtHLkG3qZgIX+BYEuHmh5echxKBc1ICax0aKjk02L
zSwxslvCSb3LhwWEk13LdCVX/uj3nLYttQPmma+k4xb4ESYlGOMxA2Dpr2P2MN5XGoASSuc8FC0o
bZJj8/KVuOTOgyi0OsmCCeFbhzX2FdXZuyMjMWYG8tEFNKtXs5luSsGnJVtF6x+F2SeCaNCGmXDZ
ehSaKU1DzixUQ/ykeLvv2u3V4Nslppg20nD5qhJUPXwpnJxMIAcsg6ozO8bG+hScGtrNoXLFrJBK
GaI3DAG5gSuG+RXc/SkWtsdwdl7iyqzgdI8iBfbn0/InQqtqwVSjmhcElPcxwzAF4F0aEWYNg4sj
odprGI6k6EJfnq15axM8HSIWRyr/HPFrPARJ51W2GNjQd61+iQcq3oLjFE8Gsoj/C4sqc6J866Bm
sKkvLMBAXovpxVsxmqsX+C1Qf3ey91AB0jMqG/O2G7Fx15UMMurCZiKim1uHeurxIIe8PbJ7hPnp
XyugCpIYBBkNMFvIcEUmwRU19HDdh7Em3RV+un9Fnu4x0tde8q5IS7dxPsyksuxZt7pRHDnky/pb
w7lHsTGr0FUlsogkHK2dD0N4nnbqVmGxHMP9dl3+DVJJNRSAU1Im2156mI0g7CF2IechSEpEgLe6
lAGJs/KMTkjTudiu6zMVeBU3U8KI2jlB/pUyH6Yk0fM1yawFcwLJ2dtaTXMQQoSYFs9+0+aZ2TRa
X19pWuIwQ3etu0bbN+J0ho1Qz1SgkYLn+65Q/Hl5tTOrQe/58BpgGJKg8weO7eetePP6UBVjIAD5
RpUuH/3Ost+4+1sXWsht4QViWRGCe+3XgH/HuBmnNrt3Pc1/iVV3B8iC/my+WSnIa023UfoDjNPY
wcSHcQXA/D5nN4TkKklRaYGVNTVTqZlAQdyik9OODvFkV94LOH0Y8SvcSBAFOLc+Pq/atxPb+VYz
gvPWTVscIGIxKFguLQMLE8ForaKC4pZqZArpkgrZTxNyGH+mLRknZcJCdJzfRCAmXpZklxHD5Drv
LsLfJYAA1lJ4scBOUrE+rnPaljtOkZI6zeNYMO/MugAPEvLTZxPhn03YMdUPsGv0/lsx/9ia0dFC
Vvcs7e289OtO4xBSydcg96Zvskd+2T2z7g+7i7CsqmYVr585YR0eDAVMa8Pr1lGoRU3XWR6Z9vvb
s7ReAoCCeFDTOztR7E79NhCeAuMWGMez9jXNqCmhQHtHto/h4TdQ/kfT3Ur2K8Msu8mQzTaBQX4F
XtZs2yaq8Jnhcn1+75jJ0fmjzQ+lN9JsrhkmXwIjmqtiPqMJXiO1sRxMicWiQIAuA1dKaGIS+I7W
nfK/3tPfVGAtnXD9pNbVUvW5Bqu6aKIB3sO0XbZJwyDfD91uUaQ3X+PvFXBnOu8bNBFWXL/Rw8ht
DnyNGsP+uuG1VN+H+ksKACRQUT6mGGgnSRCEUXJ4kJ6iofeyplOe8GyAdLCFeJRMokzuGX5q/FFU
XeEHYnCT5hoY//GT8jjQoa+EyGTuasjGnN04ZIh8mbBVsOo47yNZO5QuTxbBkqibNT5uuKFFeBsl
Mcra1zgd3p3KbN1907YQVgF+CYxNVa0p1sLqjzbQlATQUaikf++8YuWqhd/qIi+0PQQu0+sTUtSb
BH1FZw5R/n8qxrJLaA92U11TIpNvyqL5XVkGq00LuTTK0XrWkPKr9XpxJV0NZ+PfCLN+goGf3EA7
0IOtySMvCTSrTTj7PrwmnUUFPqvcLwh94HHOgafOFpngcUfkLbBfC7BmiVheXJm3PlorKbuCal9H
y8v7TyxbVZC+uX5axA6SbsuNljvXOmMJjCMxXQiMb5Q87HWdGYZGIJdHzpBS6Ykv3fzRyqMrv/Fh
NNOwa5kyxTuycvI5GnO2RlaVJOloJLFTTUxWUrEQoctk18O+GbeSkHaFcpbfLZWttBk91kZU2fTD
pul0BAYE1koOZVnY5zkDXoNhmyex9qYDCp/hVNnqe2Klgc3lj4YxcDb8Fk5kvw9krAn8ZW6daOWY
n9wef6lUbjLvOedFlvYppg5m5TFgTG3cFd8HaA63/Z8gNBF8xKpcrU9AAOoNU1vrYNQmtRlQjyZb
KcZ0HSytMwRujacnw3bi/bh2HWFI3SD5D1wskIC8bW1ITORLIqfkzyp1qRmwsvsHCpi+8ecKnkAr
2P9GTCdDz96qfIIbjKVR68QEUPdBiBFWgcPX2xd6c1JZ5uqqpCBeci3dPm8CBaNvrJaoMszfluf+
3TVZHWDBufc/cPItQyL4ODFJ8Zzecz5eCHv/kDHhJpzAtFR0mKroHML5/+QEaKBUwLJ93z2JF15n
H4vrihlQQh95HgTfJtFKueUsO9bO8KGQbBaPPG4blzJr4WjRT+zMa40NGbRZlPqcPanystF1AjaR
d0zk6solhMGntC+9G5LioOW1vv27cLDoBwLsECiTzOuanBRWmdV9jDM1qnNFFAoF3uFBaJeQwcAQ
azuyKDddVKSQ8eZHFJalubR2O3GsIqMn/CRCs0MPegjgRtr8kuMGTXzVip1y21mu6W0dfNTAO8BN
VKmyMnAYTCdSRq8zo5fzS/7UZu/XFVglC3tk7joTqIwhCebkxIKWKSqTNrJ7xuYIxGqlvQ8CDOS8
l2cJYzrr+yhfx3wyjGrCq7/0PqlJGNU3RjSa5n72zuxsc2q4OqJAPh+QyNmzLcv1KHAxy7VeTByK
jCQ9gLufigG/zRFJ5EXco7EncYJsODzQMRmRJnyuu+iNjoOWl7cjv+RJsXgOL1r0f2qKW2t7FXiv
q+0bNPKobc/4RUjrWWxSIxmmvTgq3tSJ7HayYWjvxaFZM6ZoC6ksYYwFfgh7kwkku684xAZO2U+u
yyVi0gXsvNKrsZa4tN/mkR/TX2t9gsxdGttJLsG3cLIp7aJ4MOAeNJZE0/BmtiDo02/HJfiBJvT5
CQWzQmOhZ8139jWYKUEWIi+RINWdQtZRambpqxeNGgugzjqb1u7jYcwrk1eVwMgE6AcVAe8tavqy
MXVV+S29i8COW+2z+8E9ixggNDRc/1zsyEgdymp/JGkrwDG97ObMPJS4bW74MPDVMVfrBh76NYRz
1bt9ZOS2zYzv7QU7sJKM1NykFD+SPJpyNyUVqdhgJ0xbHeq/T2Tc+LW1emA3thFBUMh7FZH90DEy
vbG2svx81exoXMt1uJkR7IYzK8iu8ewfZ7oAQsrEYanFd9R9FxGrGvvBpc1RG1zbKXY9sP7wmUIf
GFzKAg0luzCerH+DWuZ+9Yg4quCGpNYGnjxVKBiH7t6FlXjyOAgSOr/1l4JbZhxBD4M0ubasRNKJ
IPuUgvrUcoqO2LZSL+i3nf0O00UNe44K6ysqigxwY5Yec3SztTugAjYrtmGIBlOCr/qG88MTgnKw
WcFOiLC3pagtEJ6kqV+d9k0MFNlpg3vysBYss6Q0Hy4iff51RR9cStjhaNRzXwGPn21aSOFDVht0
Me21/exb2Bq73iBdlyzxNRofJvOIhtZ+UlKxR6otxTsJ3Y5YbTeDI/GKndzBlY0MsjnHdZiJrmfl
g8oa1ujUiIilNtHSKJcCj/RFVNhuMZoXaAw8lkXKM59z2R115zwB4X726ApRLx0R/BVK/gd/Q9Hv
3kAYSVYHYlCePEQgtRDLYQNRKlwgTUhi09wvHy16wh+AEB98u7+cIXEDuAFXkPAyFpI8oyQ0Oi3C
FbNAAqjbn2/jAGtNLO4V8jKcdo2xMUaN4uOC2F08d6CG8W+bXz7tZuhPZd8DVn8YPlXGvhNGNEMW
xsiKg5E4cY4l4IFp2vg60JdEEmCnAsYkuZDNSiSLKiSpdcu1HzggbF9KX5kuxP5+HZ7AxvI1g4vO
r4OK9j9tWwroJ9FkkbNwbbsNu6g1HZ5FwxU3RbmWnz2r8D4z4Ysv69h5wL29vvam1/I1VTXigSIX
VR68wTcgv1eHvuVskkxr5CakUky8CE6krpVhGzpK2RTOnvAY9oGGMxjL9PJ8x5krWLiEINK3OHWJ
RTDcyIlymAU+Jq778rgumrq+0gu6ALbKveJsbMIJTo9I6rNMkpXwl0wGDCrIPptqoxrnZghou499
sUrwxMO2KFJ8p0QG539w0lbaMDzokBD0INgv2GJ7jSp376b4BA7t1/aoaGHvO9NP/5YTF/B0yUbi
1AYEYRzuOVID+3q/aIs6pjaXEWwlBDChio2WyEFGvRUJbWKF5nUPC4kUsd8kZMneJQhYuCMrhhhS
jrfsA5x0U6/iH0AvPxCmsqtZcZ+vkMXNPOH/u32LgSHbRXJQDcOU5X9IIdE3eL7+JjqLa7sJj09s
leBv2ZDTSPPKd3Bk6QBKh+stRb0ESeAaiiZb2Rp4UdnaZlqFMtRweYLWd+u5GVnpeJ7x2nl0Wgqm
eZQbYbV1COIDDhadqg5KLDnLH9RDO0aX2j/qxOc903cWHLBVx2jgvj7JtfB4fxE2VzZVmONb4NIs
1XAHiEijaUOCRVff7S+AXs17VC4pvfaKo6ih41aGTV4utdoi0frzcTGPOazQ6/8YqC3kVCqHbv+J
FaIWPtacQgnR99OHGIuJDf0E1HE0W5wznXWBR62mkKl24cG3wHDr4dZpifJkRkWzOH+szqpGcTPr
JW0H5NAdqFgLLKfxHD4nrACX1DHlKyR1Oah++Jh9v62j07NfO9TMnPRuJ1yL4pJV3sTxG18g+VAL
W+zNZCU4+mptFRzP+IqU6r+wtr99uYag4xghtkD7sCCxU8KMriWxXmqoel25ogKnvoCwV2Ask8hP
eib8VOKkO7Haqy4xb0LZsXMJwL79p8nftaW9BsbafKtQERYq+F9CyoBnuXCaGXDP18J6Hwgaqalj
PmsIeneGI2YRXSyuwoa076dIcfnZFFE8OWId8mn/zUKkoY+XJd+CFhy0JKcb6e0kyte4WSeBo0IY
v+ssz7V8F9c4TlGeIEVFX2Tzxjc/P3JYDSQt/B5o2DlREo40p2Dd9j2Mjxf6GTiziuy37w1q3YT7
pXelSnBlixOPqkSlmJweaXOzKJ5wMf//U2cVGSYdLTiHn+9MNEgFvjleOtFrAu4zlXnSTzOFBM83
tBk1+n51TFbApX/+NSUOTBSMEJcEwVX8ua4/tN7e+RYOpnPYI1f8ju+oXj0rDvINQeDLVwtXnIni
MN1PcVEzW94zZCsDgVB2rbYY6MzUjHnI59tdXDiHybkGbJ9Ip++9JiVcYvEi4xabRErL6Ai59vMi
FVQt4AkAq4+u7brxduTKsnJYl0GwpOIwS5EiNkI0rRGvKowhq5xvslmzN9iiKSKsXvbKzKSRD/Ob
XkYGfrbYHIQOmYpvXsLBtWSqHJQkp51rn4CU0JuXtZMjkmlNk4jPLSizrA2NGbMNwZ9K8TsDLwga
GUPky2DvJwOzkOVoMG1wJ0kuUBo1WivuK+rS9HdTW83VwLpgt7qSUEsTy5I/TQtjPRYKSdDE0SQv
wsvkUao6AWmOorPhJ3x/I4E1Pgo8dEuE5JKOUXdkNpkd7MNC/WAHdG/EuRE6wTF6XUd3E+YRuFG9
SWq8DDB4TUkGLaST/n5/CELBiTG62y7SPj9V+7Tu7KRxhhFGRPgIl4LVdeCyHvcv+HWZ1YBb7sud
wD6aUPttezXtoQW6k+iPq7sznRnh4ZzjnNDG9LwQpBH10UlMcGp1DvhBkpMpTfBiw85OZ5fjGzkU
6an9byFz+jViG2t5UvOPAmlBOFuUyULX5cgg/U3snBIVBuur9iL492YH2eC9KpkxBEkVdPdghT4A
F+aTPNkssy6j/SMVfBK59MGpQ6aLL7ldJGs/bIAGhTUjNfCjbDGXJaB+QudWumUXCQkuRQut4GvV
psYPm2IBfikUJIiEyf2gghEIQEGda/ETgV0vVZyn+N8eO86cV14PBnCM2m0SmzYD+wbtvigEtRVk
ZaDBjVm5TxcdlfUYNfCnCVB5IcnVX8ZsSoJCt77FEr5QP3QG17Z1hsTs2WeFluEJfB9XfkKxMhBa
ELqZV9oKy/P8W2OVFief+LCb+4w4DCnsOE0NPStkTKlfW6dbsuTh1wpYFAFCrM95g/TmfZw6Tffj
7kFyQVCqRNdwILv8KNhPR7IvWUcHNweWOkBRLHAg0pfpKRRZQni79G8rHmFyZS9J0GyTgP1aIxlU
9ij6jYDzH59ZeX6ReyLHv43iEgsi8aLyGqAxLPz7WwdcUmMJphtFox+EbEaQM0VrnQiuoTO0CkSb
EBpl9OG7gG0fMNiNjZIYuZqTmVDNHa5nNmi7sqGyuYCIf9u63w5+5/pMBDKy3C9JPK3aNzqWfhQ2
ilaveMxigw704PJ8PBUxWrnoJRLRXke/gCJp4NbDum0mpVfW3j1UzvVgtKhEJpcZ7/naG/Ys8Ufb
rVQ5ys+azi/O4PVnDEnwKE3u3cTPd1By1jeCAczdZieyo+1KvWuALcgSa/NF6DO8W25fg5EZXJeJ
vQvSAp83bilu3w5tWiSjWazG0v64wxEXPCBDAsdqYnQ40FxPFUqIGSc09bHFcmzd+HbuWW+dHT33
VkyRfm6hHrCT0DYTr36cAoBWwcdgFpwDzLUQPW6jfl6heqU966S2P7MjXe+8hPk1qn+0zoIVHkqK
kid0yLnxj27kMmqgEr/RC6RyoLIjzzWGVYr+72qMtGfaFC4BLrPXUVnhPOKumjB7/7Uc9omZXH3D
HPrhbHivTfWnG0LBKnQWF0VVP/X6a+AfT5o4vfMESWSTQ31pZ774hdvtBPBmssoiYe1z4yT3Vi18
0Dn6QKC4vuRcku73DdRENT2KTMVn7uemmzobQ+axrmK6EeMEQghOpJrlMvyuZ9FNnOk7bxliLQ4P
TbW+e6Q7wT1/Fxr4g2wm/CzSs0nOUSlAuPW7N5GOORdpnJSQUudIAP7OPPAd/KbMOokl2gRsbnUC
F1NSJsFmxdWpw5/lNuTFssEULvXAkOSmdDZlUBCPDMaIHFa3oSzMNKrWuef1YTPSjF5kxi8HMuaM
Abi8Mhht21+uQkL8kzeVZlCoTl7vUvKDNXhvKzdKA0iXZK6mvxYY7S03ULVGt7gvgsjjXyP6F+RM
560d2cNbwE/cGc2jzldl0Dfe+hK5n4idYsyZBHdjt6EbdD/ZGAB6Jqj7GZLzYJttYL+cjhnd3sp1
3UADePJkeRhBaZGfFIs9tKmS83z9zhiDgMZ2K0I99RDqrNP8FMNW6fD2+IzASpsi0VttB+wxYcBH
DjaYkTiEYBIMga9Rttmnbj7kBw8lQBJbi+EgZNynC2NfbN/CnwnIOGIXsYxNQwkK4NyXWAhKJY/7
bUKPVELFf2rTvWQ+Fy8JuPqexkBgcIqXb24RX7Y86FO5xqTfnVdsxFZxhNluBedBeEyoucFLPwq1
Z3ghBDct8q5EZNh/WRT7lg9Qx7T1djUFiS0od8DWSlrSo2BD/RnZNdnnaFjCYMzJruqHHLaW3rLB
5Gt9I7kKD0ifQ92Ej5CBSJD82sblVAg1rJgATYXBQPX7jaqL7pHGWP6qddbkItVI+o14I4urwBNm
/+xZ4oqT/bzuRuqd6xijG/4P6WVS5FwE/o7sbc5b/Vp4fPfTokE6/OT5LwWgIwQ/OiGVqyO9VXwR
CjJ5FV7maqbG2IS/QJIA8Rq1w0mZGw9L0g0klYSMXFP5c5GCM/bFJ+0Zip7YGikPPp6HivAqcP59
WMF8BG1VJpK3gH09WpPR7iF4qC1ZDugQ2ZjyB6HHX+ZZ4LPJwcbrD4/DzEEbHqFMK9Y2bNPL2Kxw
AUevGkyuiuUyMrSZmvVzdnjLekctFZVp/lO9TVEc78t4AK99pGw+iQmyR+LIT70Epo4qbYYr85QB
80Fej+1KYSa9gkXkDC5iDYMvI3llGyHq5Gqi3Gh9nm+8vPtxB1OmyE8vSIUUgwQEIYJmurBUJT/b
kYq1srFNyAg/nHBQkJxq6Oi2unVaSoQ6g5CeMoKrzPzbF5AKkVJS6hf3CZvK5J1WWoDKZ7bNDnGC
+5IGqnTshS9gDEwwWiUYYsb0Apm1BUNgGsjfWeBQ+v/yGLOU2tsjk2pIxXfM+Ab9HGWMwq+ZNoky
deks5A5RAUTgwqxwn3rwu/YUypgscrr14m0w8Wx+WvgfKiF/9dGcND+XrMDlRg9CgZrYHgPBlXmq
3yVJGddohhBCSeXj0APVdhMoOmcT8xcWnlSHCz2KuErcw19MFd10zDcKhCxg+PRgqq8H7bFxFINF
arVd2PtLpSQoOMJ1rmmtaopF7af0vPU4ufHgBr3giV/Kn99pJlRB6DALftAOrB/JApjw5Y9kmjui
CpcS5zWn2sWrGukUCZcOVbrZb951gEc7xe7f3DmkPKT9nsonFu1XcHQsOtFpe06Z8L5tu7ngEpak
2CFceM9lDi1BaaphI0aGURFXPlzywf6MCemB2doxE2Cob1+m313lALflMsm+CMZRydtlY7Ln79+2
o/2QAbF0HBhj+45iHWgwx9YVCExmFK3S4MnQVOko7ZecjB1FfUL7tRRsLA1W35xYHffwBN5gKaUB
+kz1FCyu4tYV2ki9nwClpB5V+1BrA3yK48BYVUrn9QOYH2A0euOCO8WlBAuipXsos06CgL0VKjy5
xuNa6lziTwnrxcxA++gSrK0Qk0lkjXHEHBycwfDO/8gzaxkmpTg0z/zASoPNiKFbC2rutaU6tHIn
8gHGVQ9Qiyu60jLrKYQVl8KkflcKntWf/BlVFhpdvfkr4Vk5xIsHda4aj5BO+qldS0WF4oA+Yb2R
DFd7lxrkrShO8cRhH/k44+/FFopyFPmXzXJf3wD+tsTNFVpJ8WdmsQKN1sN1/Ff5dDINNFlehIv+
5ZG0awY+J2nvlhjHOWliyd7JzYDfBlYItg0kXIWV6Ifp7ZMTjNRScRN8j2V9cmlmglTQxKln1WXC
MugIezpGhW4TLBcT9cPPkMEpnyfnx49fuEET/341lGB9kxlyQ3Wl6ckaYAYPTo3nfCJJeIDOtVwC
MRYOwsOe1Lqq1RoXdBjRMzO4uUTPEzIIuALNlHPMvgf/umyUrzDXLIOWXKWaMGPvg09UBaoxm79O
RcfFj2cPGR4lJb6h8Zn+wh4MaYGkZcDDAZK912sL7b4AbRAi5r2JlknUQqGQazcMcEP6yjrPnCR0
hBF4sa+nmKG8oao+wuLpqcg91PoxZMCsfy2317vx62jKGIgqPHJk4Dh7rJG+SG0kUzRXScsJD5Gz
V+6D2wSFPx/74KSqpOPZkcDWAxcmTTESLHwxwdNwY8RBFQjm7+i14cvG5MAa6S5NwBo4W0FNVv9n
cZHod6pbFJT33vKhnml6y3BFZABJmH55NInZGtvE4ekBlJfmhfpNNsJXRakhueb4n4DfKdYXOLlL
hvwanjc+NskjELB5jNtFf6j3JI5FU3OCa0ggYwQLud0yJAGLts4IQhTxVgO4iQ6hFk38+jfPf3An
bNrdtrOOVDlhv+RiQFGl+Kqin22iWdHXFP0C708I1XCVBifSUkGoCAEP7jz9ZHVS4VpBPSTMNRze
a7Za5YozxEdBEqNFiRLCN3llNGBQT0/B3Kxt6nLdX4i8I6xbZ1wXW/N2E8XUWsZTZ8mu6z8NSVTJ
1W8hCdZ+3OCcbm7IumyvexoGbSwD9MdwEeZj9g4y4VtxnxrCoYue/edNiVYSUJSz/n2vcVyBLG2C
dx2xGFaCU23VDFj/Ht6ppl9uoLPlcOYlTFUrhFarpSIIbm5QlAWVb9omJ8T+3K4sszga7qy4Avp6
wH+YD4HRBtveGNtpDuWCqlZSaEzegPLnE6hh8lNDl6DrM6z0gFmVgQ4g2rPi0tx3SiuQNwwj9VBv
RSpwBTnbUZGhMJ4vWGEsHVLwzEyCcH2d9HtrYri8g1r61bzNw96AYAHlZYKNIpCCS/X1mnL1Zfum
EmreqE1/s77M+De5WQ5qy6zMD90KaZyF4LW4Uu8ivkOkDpHT+YnpMozR3nEcgPsfsI0xn9BxVFuv
ytIYDX9X8xClhFMjovjWKm2ti5jHeyZlr5vwjrn2CghDn7iLHR+hX1LVZ6lZp58k5Ow/7KUQkTYo
rtuzU4JDIBWlPceQ43wai0204Nz2b3qkPkOCgJrdSg5AMENfOCeB6MR4T+i0Vb8s0OPZNwtaqgGL
qENydvEYQVrB9/EbkSldlpcNLkhZ3EnUfErmN3/5ZqcrOTE/izt9ckkta2YgMMnYFgt/YFo1TFrK
ORDymqBLs+8qXHu4SY9KJDZyKW/LICTFYJbO7VGSm9qXH6uX2J72HNiCm0/dv3qpwQX/Djrhvj5Z
k4ikGz2p+hE6KDWta9EykMm3os8kPW4mIwq7grLEi4UcTfQtVPWO71arEgMHVRAV4TiP03vDfkjG
U3Um+unbVhhVQVUd1/1fndlkc6PghuUZYEDys3Zupw022DaeSVK6wAxiz4/qOx2pLVxJBB47b8rQ
KzU/YOzUvaUu7eKXqk095jrAMd4VOW9aQnxuF1V5/wqD3vbVhNq1cYe2K0LVL4Fispv3xarqSlC/
pSgfubgRyUeqBabpJbqQQsSE4pLIDD5F6kRg233arf6mH7oSo8m6fhcc12flD2DXPuKqEBdbnT2e
5rOik9HXjuwpd0Pj43edDLtjHN4kgRhzPu38xroOajv2v7MMT1S85YjfcsjhDJOtOTOZyW+6gOD+
PmkmQWH6pbm8kcYepmPqpjK18FvumkTB++9V3gVqsnQPxobRrr2Ef1zhzU/Yz6fXR6UyDClbFNrG
jkLwup0eC4g3qC50Yw1B1l/NILImAzr4Qo7C69dtYIy/VE46BT8dJU+Y1lhG1jW72YgBua8QIIw+
+eN0hCJkO+Om/+yhIpkL/xJdXF+nC6Xg8YsGmkup+UwFBJN/nLuBFkyQfKOBiabFt5w2KsZSiX7n
FHC9HbJW4eil+TNHh0ABhBVkyJdZW8kEt+KnmURb3fjSLrMjqXjt6pvvgAt12jE44nSiLT+GvrfP
+Vs5iKDcgWdZO6+BWCHge0TMSotRREu1jL7YWZyCi8hGCeQ23tMCrogOvpgjOFvmFPkFCRzLmLUA
tpjqY37brgknhXmtjoMYUIl9bBl9BxJglozWoPabWazxkYnQSsUz/jLuPs5tRtdKqaRNreaKhn0E
yU44DJcaPKSo47scYMOoDr/m+YhvHghe5p0ypt9dl21aZcDo8Zs5G2Yz69oylkKkNm/xPHjJFW1o
w0pw5q1SRcq5py/KlyIz3rY8Tg+Wigt10srlSedbssNrutQV7ZZB/JicjvudB+jTArZAuQc96Rsb
Ygrfi786vNB9Og9ZD1lfyJ/3C1tZqq3rK/mEAEqy27e7N0W3TMq6ZPo1KakiQEjAXW3r6Fu5HLtp
WYOOFVzD5UIFkKxViaNljrchUVECBZgXH1bflQQHuKSYWnitvlfglL80V75iOX3t4IA9f3lhpEKb
lr+VUFoS+yGkGt/3EFywtYKH5RkFymJWIYZ2FHu/ZYTGekl4D5JhJYfNik9yHFHL91OuGTI7iOlr
SUUi7yF4xAkZ7b7mRQPU9GL/j6xUeNsXpROYFMTVlyWi6RVhJTEGnX7xXpoc72izK0COmnpNdfTi
ogl74tR+IvubfdGVsBMzwiJk7vWF/dLBMMjXIreubJVxKKMImfX34iPB3mnAUPpbdwdLZM1yMWmT
EtH1JyLI41Gcn7toJtqjHLctf9j3Q+qxzAX3Xe0oCE2L0MDERS26AGIoY62d/2PbVuow6Ue7LXLK
L0y2P4NNIOMlJnv4z/jnZua/mcScnInlIwIXF40faJJsQwdJ+sJkzT8Ws7z1ku2c58k3v7186EZH
3klHXeg2NGpB3SJh3sd9RtiQ39zXWFYF1+2h6Zdtv1guB/bMnUPMn2dp1OQFn1MGfqD7g3+bi1qw
/F7si7GHkbKPqlnniGbathGQLUxee44jW56uVhZ8AzyR9udxJX16S83/a3P78ATo7yIvxzc02OgM
HBH1jD8qsV9QKmCF/uBHcJ7+eYJ5ife1LsiyAN4cfsJxGjSOYpTXlMA4EnPJwIs0aSh7ZUV14V6v
wuQraeS9jWJzOWvp4oqhmLG1WK/WLF6fJMhDfQ07QuXUMUDymtqE4fiJ4kNWpowBlMGc86YKmwlx
sKF3ZPK9G8hz3i9bQQmijLNTvjVqUPEMknTnhdq+6uRIyk7tkAO1yU1CFpUXU41knd4CNaAg88jv
0z7edoP4Gbkj6OL/AwPCVZ1UpsDYgmt2r4whTPOEErVnU2fdetKsS8cuyiK1urlhRi0yglpTZTws
OAl2k8svxH5AW5IMBsS62TgsKZtvId3hVQKzpot/qxE9xqWeT6BRui9rnkUiu05JvdxQTaLQBNKL
OPdYsgmqqnjBiaepVOn+84aeW9sfzPaqsKbmQlV4vc2QjQIee7LzzM2Y6RE1t3qfOcYP1A7xAhTb
21Vgjzzel3qWNliRGN+Wy0iBmE7N9eX08K9YE4kvSxLDoqM2wWrbibqQ+qWuIm6cMPcReoqMMCU/
RO61n7EfmVy2W16Tk9NtBNXxST3fxYIDjslsbyjx5rwH+/X9SpUWrsbVkZ4KLe+j7/WFDicsPXDq
9wY3RbOfNMrxstD5m/bPk/Hc5AgJOG8l1rlX5zB3pi+WorZHApQ5bfIMR/5UfVY5qiZoYIoVOgTT
EafHtTI1UJkpeTfKWpExqzHKnxWvDHQLcUAsNclIYp1Yba/2qI0e0Dr9kXszzOFhzxK+oLBafAb+
oxYhLkUVbXgtXYNev05A7E2mabgmG/WQ/M7kUVzh5qaA3+IFZjlfSitrgVgNfXmG4T5e6ZrZdh2a
8tFpChOB7gQc9V0DGScYgjbkyUD3oSJlN5OBflOoNYXWyzq21ZOeuxEGMdqoAxoWYT9NqZOJ9rQj
ql6ZpbHVe6nr98nFbEVub+Zlq+ttU07SCeSblC4hEAOPGcaI9llP8VUE82fvbeyNG3VW558v6+vO
Ihvj2iFlwdBgu4OawSiY8LfIjOQf5vu5jQPBfCx8iq+cj29a/ROqjRfawIX6Fq8D1jS606KCMGk0
zRWRc7fMtri7w7snhaEkcMn4up9qauv35deAwi4F0EAA4qhfBl26urRFMtDhAiGgDS7nDX3xXvSk
UdCPshfqE1ajIFtljZF1nL40mFtCgmZNObz/LD84ADvQJx49f0Br4UimPdq6sAh/xxHc0s+QDoZZ
whLhu/ByEyk6mwxHF7BSEYGI917Wi9dqxgmU0SsqmyN38+kEjzWZh85cJknqWR1aMeSGtk17Tbxf
kLJ0vCCc2XocH9Ekp3zL0GytFauVnTqt4vL5fUcwwI9COIqKdYEcg1rnmKEch1eMqT4OSNm0kwXX
RL/lQn3QAcSOaTQT/QRWyYXqnMS9Tkwb4lrSAPOS6xGm7yZTD9wLLhYCKqNKjbsOelA2E2Xv3C8B
9/itpVGA7eeMJzhTXiE0zJyDGGmZPE2z5XQK0UjCbDshGQT/gfEayScwRIWR4bpW8YLej95WOeAG
HjMvWcODka4eO56+0QblprJln3V3jrixpH4PyhsQnVRRH1RIcjuu10F+tIEhxyHWkOsIDZQTBLZM
ks4uzttHwLBx/VPMXazu/+JZdkApPney6pcQ9bY/WZlAuhpK82dwrVfmuKolkg5iL1ZX6HgiLRdZ
gXkuJWaN5clgINW86rU/PAsDe2CjjEPHmMxI8hqS9/IhsgQq3dlidWw7QaFDk9Q+6sPw94441SRW
PNhGfV8v2OeZvlSajrHRyUY8QxccZj1ykDkSsMueLN2NfXbul395JJl3mh8aIodU4oy7WA+5ftlo
9zLccREzzsqSR57/4kkV5zoZoPWj5hjh9XrvmHDQdXBy4fOodji9FbQ1JDXPYlRTMCtU84RoRd81
+iY6zUhDHK6/YL/3I9z56tQSu0y58WbIZVTm/mQxFoLhnmejh1ynURZ8d4bIH6yZ3pEfM9VU69kJ
sW+DREUhwPSGmEHzCrpZZoH+xEX3YgPvhc+ZV9Nt4qHf/B+JP9XoL0PlokHcWbui3wLVaRcg2pLu
OE2Pd+qoQ8B2qzXuAi9QXbCYLxb6RgLInQzZLPOOlDAosn1Yp/dPRK3lxUIMvMmKQ5G8vYnyK14p
5fhuuhxABkMMpdRUZUXT3xgvKm+boYdl1aVa/K0bYiLb/DhcOV250dCS9alyRmDTM1VFtanYAVgO
K46onCvol8ayIaLo72ZvjGxYU0rVKduUH6HuYoM/40h+9w0DtCtdBTzujzoQsvuE4rWBU6997til
SiiQ6gc429XqwdoEGMzY8b9x1kO7zKaPKGcZdaHk53bXMrTVtnYx3EJFMdUKsUcrZ/1LFKVFHBLP
4IKs4J5Mm/00pvApNhxPFbFFAlMqnWvVgEGH5SAPE5/3J2O0UnyGd1iaM0XhV3BCy0vxV/EosCY3
dwvIgbwQibteyKqyMUky+PFi/18+tnicTH2UAW/PudH+7johQVNRVrcwrl9Fszh8zMBK/Eab0SLo
0MjTLkJ3ggGEnSU3HhfFNuHmJox+HKA5aGtv2mtttFukpLn+dyc+xBNylgJyuln+3tcZwP4nU1oM
QqNLEed3GpLbVKw1TByWkB7r5LJZLWVrBkNUSXfmNwwRqGt1UCumpc47Z6FH7j1hrfFqPCZ9CpHA
7wBpNY02H3GuJ1BNPCnrj9egiTzYRgubT325r7CVpHnrYwotAjADdBPwwdstqNokm7wjE1AfnnMm
+Gte2eNxBFKSxMLVb52EFT3kWTWPLXSruTh0L3jHO/gvsgs6aTqnTK96MkS6zmVm3NBW8iM0hN4E
THEH0amR/VsAI8BU0QvH0QYfMc8CunKeKFHUOtqziHIoOfg7R0gb+pDYor+69ehmrKDAMg0TmTZR
zRdct2njeuu09F8Em3HuN0mmOikA+gxNXnGD9cX5KtNbbTwK0qCmgvD83waxEpt8VFVVHBM+92LP
X7cMKvBat+WuBeyqN/VwUHB3bpb9FC33Jn/1dyUP5Bs9UhISjFXl4G1kz7ghdSGxFX+ik5aqes6V
NWnLGilUfigvGgkR9jNFezwxcRM1SuMLxPDPHk4kPWvYSYmr/QWJ936xFbmv2vtFok4Uj46Ox0L+
AiujPdQbKC0LUNp4XwWLTdZJSfKm1MMuUC9AvXEGNJe+ujaEAve/i2TRXEkWbhStJdojQ/liloVo
paSz6NlS9XtAGdp3evh9SBzZLun2SBSab+A9Vlw6IEeqXOSj9Krm4iSJ7p96zJnR4DGO53kGeyRw
8WZxhosIKuCJN6An1/f3X/pNcl9apHXBuqw4ray7hW1AI7LIlx44e24fNtjFk9CIjHC4Mh7GvQ0E
yCaFNTZfmcjrBE1ZBuC+Gdy9IxY3tcDiTWc3+sbQ3iUZGOcrpeWc5hLuh8M9T9Gj+5vRJQOIiPc/
94wTHgrZa83ZfjPq2dGq6ORMeXFBjsh1fdjwJiBd7seVs3DBLAki08NmZJw7plP9Y0V5FTGVroPv
jY8tlnV3o8X9+M31UmPowqZohb6aXyS3azu/uKA1hPeMCpzX1XGBQH3Hi/C9GFdJldxUD9K/Bpin
5wMIi3s1cUot0rncQS4WdBgXHF2jB4wofniKUsVpz9/SeCgm8+dTHP3cn0kCS6ABbdVyhsXqmwgW
Zg56u9jn7h5rnkyiNceajMZnyiuNnRqFI4C54mDZi+PExki5xIIPWcjJdj6snRU77tkRuqtS4QFO
p6u++uqGv9PHUqhXx2xqGhh+4XK4H/gPArW+leLGc+5My+NVmjUCjzx0cfM3JiWklqiZSr2g2kYJ
PuhCFRbSRtla1+i4BWyo8MnbfOsWWkSyy3NxUQ7dMVJBW9ewL3r/sShI4idln/H2nE9BiO54e0F+
RdH2Lo4rtgsf7Y8fBWvabpOCv9FUkf2NG6DdTM0MyXOb4S8YiuGBKLOAqE6BsyCcF9+Zph5NeAJM
9ozC2OMjr9u9MT8xUteR/b/STOwTAKCAvjuMnK0HHiPpmpWPz9sv3BQ3cEztDwxZY1YFrk+c5Cur
BsYnq46TgLvvGMMGnXLFMJhr91UByL9aQ6/IuIVllr0QYKRrKzoMJNwr0LTWR1XXdof50uw3ey2F
yUBI8J2OzD5dzUL7lwdMhFzjguamFNkq4U9xcdU2thLbfJuzN+gBbvTFEhTY29bkOaxITLmOQ/6K
wvfA/gisGC5NE93QKRx9yrnqUpGsuLCuZ9J2+PE1sr4A5pxsh58RX76+hv304wAD5xvYHOwRLIXn
laAT+qW7zPb+QpkJ9XP2kvznZDJt7ZhYHj4ADt+8Q9PKtPIiw82OAJZHpPJorp09qV28yFy6eLoz
sLx9SN2GH9kGt57hpcrzgU5ARbOO5Taaitc137EPVzOqWP5uypczly2GtmJrTAYjW2MGp1vI+OOc
h/Yl4/WrPNwB7TSqffeosV+rkMSIvzMTEvHO3LZS6FCv2J2OrRc2y0/KsGXbPkOnmK//O1dMA/xC
Uhg94heZ9UL7ylNLUmMHLBgmeCb53op6F5ReoSZVoyNvy+qWk47CMI1bKzTcGVx0jfoOJxwjZzy+
10jN0Moej9HOD560UsFTteDvVul+reMRWsWqUcozggblYf+ZhS9fCoy2UMv1QcKYUUX17alglnI9
0G3cw1ks+LrqVL4dwd3v9lWGG2a7dtKYeXahOh/f4Q5aL2b2zfsKwYMG88AHPwuzV8nKuinEETG5
z6aFEz1S6bt7lgPmBEbGlYOceHLcnDjfTte5l363ZI3DXChUikuYV1OI+OzUcej5ioXMKzUdrxi5
8ifIWwzOWAHFdQGs5rJbGbh7rD4cJY4m0f4v7vKK5bBQgo8poHzRM1I/17TTQPbQWZgEUTzO8Bhm
NADtbjbftKT5+t/nNUL49V69CuMpsQgj5zVA/xadzX+t8CtpDsMlNiJo8gFuE/dCEi4IIvmrRuGh
HwgMEVtpQHsWtM1wruVRCg18I3G9YAmdx1EeaTZwPow+GeNJlBijssvo0AD+Wjx1jsCcOw+cDQc6
lPV/+6soqazW1iTAu+dtfje/JFra3xaLc3aJ0pgsgC82MmBpz8oFBSJC8ey60Q3YyXk7fuu0us5E
YYL43CFhSMqu70JDUEOdOJ2OAj2xnY8wSPxKIHJcm00RhMTr+MKwYSDgl+gcySrDmkVIlaYwQ2CI
F6ZApvn90clO8jsPrt6Te+yCtmFF3DQbtWqVP7fnnL28OjwIbFdtAjoAAZP4yBj3tRAd2xXL0rfq
T4ZktLSNGCwVRo4ZTHRiAU2zGkWX1gvvha+ke4O/rYYhMaynfFSD68WnHBdGa9z4M1ca9cPsrDfw
uL9pLxEXsQqbd093LYJkgSUakjzPOgJQWd8WTTWpBYxv+QwweQahwq6Eobp1EDNI+QRO0kPZJODA
BHpuU1hmLbLmeyLvfmp1Db2vasUxgVNQNBA0bqATJsZsnYsIS0/xiQ+Z3mlbbeu9PuoJwWcQTzip
0mivADOjJr8gUJYC2V6blNSAMjXzOqa3t5QK6paIsWwzNa8Dv2NWHRg4JDaYISHBatl30ye4vE+R
TU+UtUe6tDNq1rJekz9WreDzmv11b8mN3LiMaFS6f+3izGB4ZyPokRp3mb5KzF8jKDNUFOMWmH7p
7+u3Gx+M/sXtEu5nQG1IQp1goxn+3z61FqMbVUABDHVP1lJ/oSlWHqkn+jOR8zRRnYu+u4VyhlU1
ItOHSc4/y5cmUMqqesXyxJIlE/t9WB8EADOWJuQ2IFEKYkQgiFKdGBgYTcos0vUvehXe1FiOJgG6
tC3DRSWiVrmS0morZ4wTBgX1oxFLPqEPP6i0eLt/cr5XAsstgpZH9RqqU8Pq2JHSTo8ConIb6qnU
lIAyxemG81uhvus69bBEBg0VTEuxBwc5afMZHs/mdVrG+VUYSzhF3wCJ2AiYqzKFUblELFItUmM2
DA/4EX6I0mIgLqNIGgiyn+U1V40cV/TcmqvDHw7VS6+AL4W8VTm2BZcwOVn08jP4ssD7umz5g2Oa
uCt5xId2BVbsTdBS41xuvZHvVCH5DWfEku1tJNN6QGX/5Pqs41x7seCh2Vu9OlTOyUozuIHRZ+sS
I1zcnmKDbN6jckMMfGNrkMFflTIwkpqyhJ7V91B09k3Nq6oc3URq2nYqsOhJZCM3kskyCeKHsmL+
DNfuT9DR5cLet9MAdj8SVzlu+8z/PApyxDomUz7tzWjEoeOE/QLOV4nwnylQFVd0qGjJlMBe7mxZ
azp6GvGfxkROk3lu7cqzLWdw+K9b+zFBxHkvmY/BFWHhY8ZuPVMDuclHAvCsYlz/SMkGz6u3W7jf
IouNLIKjxPkOQSgG/M8n5fmMqSacyma8dWSC+E2kDI0ZU4GXJ5DgSg97wuD9/eJ33iCU0LZ6yuMf
o6X0XjeOoruys4MW0R/vUOINV+tZF4fF6V28SWaFIejrkVn2PEX8OFEPKsqxuyI1XyvEdkofZu4+
wp0IvlBnLN75HuW9HbgLiRfm2otoS287hQwufHMN6tw+siAGVM+bBjWQju4OpA4Eoh8QP6prizR2
RFvPqnQ724MJ8QJ047Qh9PMgCA97K/IvQlYJcca0YkOdvxm2PREA/PEOrlu4pI/29fJVJu0f5af1
TW1JwrHwY9WE9s5+RVFAu2RPvHElV+KdObMAIRThGU3BFvqeELD11kRowcw9jWTYPlxF8MgEQK0p
zLJ9zBzmkD4/80tYYWzIWtxrLsIGD1ZNCSnAJ6nGK+axibeLWHzrFVtUawFjzyG4omZp2G6eeJux
m1LRD4B5poWHxCB7xDavko2JK+qJ3Jzy5t/67p3L6HU/vmMmqzUN8HKvfYYOdcBg/W1qFQItFRQ4
BF4nslxP5Nrmf/dmc2ZP9/+NMIPEsGdCzPcOstfZ0e7yOga7xTBKpIZHKNzFaBelHJ/kPoW3L9Iy
ERRYtqIRtlM0DjwXgC0dyqs+a2/YX3YTsuE6N2U9oMm7kQ5UUNtZxqIG4WuXrGUk2mZLpqwP2ybP
cJb3y1nrfmUMXDjK8WjUA8QhsMPEdPjOmMfvYcAhK4jgxK1bUmZ5Y5VXTV1m0xgku4Xzo8wTwwkI
sFftqAZ9cp+LFHBY6aHEVLlGMd6elF3RtVPtxX6vXMf8uqXQX4rOmTX7KVPCD+EnI9ia/+LDmD52
rsoGihczfCtUHgV7lMmN5wxK7nChfdrbgL65czooZoOhvbRT0Qb+ZqgYH/b2oxhzCwXISibS+IOe
M0zafn7pFN73LT4+SiZH1Ato5JPkL2Y1egV+AfeBS9Sx62P9g+cWmtx8CLi8eo1Ek9D8d4o9GYhm
1fJpY43TzVREuIdFN/G393KSjvFY5Tn+SILeNEY+cbR1OULOeuaHjIXlImTe1SvqAuy1KfSTHJ5W
W2Q4rhIvOk4/rzSKnYvc4PSoR4nU0C9gZhyyC/3tRIsjATbSYoejDlrFoTl03Mndkvd3igpBvRgi
jtDrYB62d/8seay8MXrXCZNZGteUr7CP1ohEEBqUI8VBXwapp8vK1G2NdAdrnyPwzOXoJqgDHl+8
Jz/M26DKhI8WvUyl+ikdKNpEXJhasw/WyxMnp3BIjqdj8bvqRH/4qyGsA57Mz4J+eTfgfNRkLKmf
cFDgJTNhMtNQt07mCfqMSj8uDTJZ/llTC89weoaEEhyfjq2YdXBytICcGTwSZ7sYrEYkvpJs7GsP
ItdFOptodPcGcedcSUCfqAsbCcWiIXJ0VqdF9Ap8oAJgWt6I64SAQdfdVxgOT/umKB7NUx5C6nPZ
8f+U2J4W7JFTI7AE9bJeCV53ADTLybAvMfDF2LB69iWVqKN/4iJjWfcEc3t8I/tNgMYrhQwNQkVb
KpQDN5BN2ZbHITbadkd0KcQj2RHkc38tkCejvEMpmwgilH5zaShRVG0l1kebizBLLmB8uRwimOE3
uPoLoTsIvo2+VcL2hpw9XZQDldTnUNPlQj1wO3mBsuKNAKsL4Cbr3SJVc1hK/yY7qgIoAW0Wke/j
nEgEs4v3BqfIzLeQrY72dohgIw27UXn31X8FvT2XFU+g3fPZvdbFUTldTrAbXxz8ZDgrIDSzkyhC
aIi4+Og491TyTsOvBY0GLnLMKI80zoamvb+ynPHGwK9cgp6BXUakHscPlQPLQN1NZWsjVrQk9f2I
xUhQEW7YtfWc0XpBkKb5KLHzYtwtnRUlc92hvknuaUKwnY9WFxO6v5aUgqwO2jQepP3MXVbF1fMP
5PZeynYNP0euGcbdnpZCbxVMSCKG4ssLPn0oOuPOkq6YnCL3YJs9SvINBaQlXJERK2ZgLs/4lvH7
n4ypOzSwDt01jfNjJnjR3bh4WzrUVX3nutuGqCnbWZzmSbVmCPT/oQI+0CFEFP7OYUtT3WPwUo6Y
VS2XXOG6K8ZnWjrO6sVvQL13bHC3rhXeNFeom5C+nXHam+Mba8al6ZGhXae55uv6f64uNpIxqeig
ZfhS3XoJxj0dgKV5M+QFpFmdE9HqEVmhD0PMY4iuT3vMbCUGWClZrUH0oP5QR/hlNzNw5bY4c4cd
mL2MhOBFkbmj6fM+JOJ9df44CqXrUKBdNmfA91Cd28ZpxakL63Nx6Xzh621hyvHSotKTtPmwapKo
IxBT4KDQUvBXaMbBISSxlwym8ZRQn8TDCkCwn1orn1tpDJcIBe4tXSbpNRb9/F43W6dur4420l0D
P5+rtEO5jzzrEdAz95pnJZ4zimpIsKyK1en8SJtPohWciJKk5PVqBZXT4CV5Jucrb4R7nYdq9AD4
qrYy0ylyYOppQHvY0uF3yzfna2OVAMNTUGRmbBdtXAgCd3ylnG6LtCe/FvI+1de6ulNWkYY74mHH
STUnmHa6HssFbwN2lOA1cqxh2d+InL8pd4Y8Y+Hx9/BBv0aIu1445qoG3MWMUpaS1jyTm+SyCMqa
LlxV3F2ZiaSM4s2q4SxDm2iw/JPotEdPPNQEaSMVDdwbTtM1I5N2BuKJTqYy0hqMLhiVlHhy1wYk
DEjgBnpLgfR1qg2VS77CbyQ8QbZeN+YRTggZGlsuq93ed/X9oo9VzpHIO6d/mijnrB8Ay2FOjwWk
Yon90vlsKHvi/cXbKPMvl/D8y/kFempvQ++gKfGmkW9eFc7CGRMG48UxFojSeikvDmzBjK1Hbv0m
pgPV92EQWUtGT3Ozs+56UAQLW5UA4Qh+Kir+JELSdzwWtkT+PwdJ/fbc9DsH0sOBKFL8PE6kbW9X
AF+orNCUUhVoA2QuN6IG3hOzout0X1M7y5ZvMJOwMZHa/ZahLkm7Zq4WS+FK8wCXxhp09EQkmfIt
1Zy+pdSwAhcuqPo46THp4kAFd8izeyz7UGFrHrxEasmJ9ZC3OUuJp8PuSZrYGBfHHGZMQpNNTxiP
tFn2s/sOhZvouhQsgHm1rwfGxV7uq/Odg0ocvQXLIdzZfieI/8qpYLHkWzKknCvGlMsl6ng3LdM2
Zk1OQ8jPtnHGRk7GpT6IrWL1LkCN5vSkWM+qI/qCuk2Tgh37H32jOgQUTvyfIY8hwYH9gki3XqiZ
l+dTjdR/WbWY8C4CPqZ/IlK/Xj65Zk8eo5jtqkbLW24K1zT+frbsESDK2cvgamddoOTGumpb0L5T
OzKFv1XtC3nD361FHowJ0O7RLP0Fv7MDBBtOr+X4XQo+EiajyKzLI9ASc9IvWONfmiP4Lt9yxhi2
bJyuEdjq2yIMpk3c/MP1/BKJGmlpJaLFcyPDC90/VFuXfwMb7nTBp3heGl1CftY0Nug8vSw1OWP9
1f61LRmLEMc0rNCxpGQ/oOetMUJ+NfzncCD9tfuCbJazRKa0amsKt5df7ljtUmZU8b5G0zm3se6Z
Ns306s+PCWiX5q0tCtGMK6qKbVdaGTFTiznOWmR+AI8KeOJTXg2J8GyFXyXbHSPSxOSxUd4OhQ9p
0tvDVFs93WMYQpli/rKzGeMPUVzhkpLUEl39z8mGHf/0HcRcf1wtG7Ji1eRNH/+93vEuWmBWP3wM
S4dshYQrx70sjiZ+ouLJbp6x/4FdfCuBAUW6tao9dzsPEKyNW+eo24hKdx0kQavWFw0CBLNIBHOa
f9qmzyynWtQN57zTv+rSolsNx3yDXE6knVIDfdvNcGi7r6EZMOYBgTIew84ko+JYa28TFkGymw1A
UPb2r2VDSiRrmQ+AchN8obxGEki2EEASa9akvgi+dPHeujUc/NZQJXALN/nSYaLotM/jXAf6lspq
emUUyGUaNdKN3YSXw3DLarFhwQZtcW3IG0qeHyU7xF0uN/kq6+ke6h46BbqXl62C4S+SKzYEDfRF
x0d8Ajd/P/kkSD3TPlg8a9aIfFIDldRd3ChA7Ui+s6uU6Car+8Dgf5Fpt6e4JMSNfiOTebgPKHo3
Qkfb1GxU5o45D1A97JnaE566LcevlYZFLR8Vgs6R1HlyYOqfn0Ayt1fstcwmtMNYU0WBEY0UV4gU
7fn3HC3TInzXKm0AwQLiEq2EMtSZ8/SHaKuVDIjM1X8edTwG1dFveS5amvtkLhQOXBRr2jPoB4za
jYkguDOrNPWnPpcrM3lL8j/7m43P6g9178iTZkCAk38zR5R17dfeGb8uw5BM4wnyTjCwi5LkJw2q
ePdzb/WNHIsa4wKpjkM+MrzhLqecNaGzd95Ce6R4lqorL3l4IaAja6uW8u6xxg4afGdIHwUKZJxh
XBmdDK4O+88LSUGAQCpH8CXiV4zuvfbZDuQWU5dn+5udDxKA3GjBAGrfMgzZGdtXH/tsI6gO7E1U
dTN5Ez8KTepZzKX5zbnKd0Ls4lKa6kUlKpKX00Wl4zLAs8tNMU6pAqTAJHjWsLPURMXv2N6JK/TC
5tARcVt/RNlz4eYlUVH6yKaI2F9OQ5/56tZ7+RT4eUShfimTMF33pdwLDZFc5ZcciAegWBAkhCDn
1XvqzWWedI8j1EDg0cwUFEJyBye5nguWRYAmbGKWf+JJIU2jphKKgTNwMWpgNzVblD4G4K43VoR0
lPq7ueyNyQfYpM+NZvJ1IaKvzzUqOaT0tSDNDP/0retax9zkWMTMGWHdbo92cvZGOokpIxZunXSK
1stV5ThitOo6/OGU4paj9FxwJkFsfzg57Ciz2cbaeK/th3plXG57j70R3jNjHgR3Aq5sQkq/En0q
VPqbc8yPhSET+Q/pDKG831xYkBPjKHGGaXo/YqlyUKSCqsKNCj4exTZStdCt09vUlSDw/J/RTyjm
oh6XE0yYuXOaoHTyRdeh2h78x2EA6Eoa109NW9TBRqyHcxb4M83nzm3jWSilxUeHXSmGXDWABNAx
hgyrwNyrYy3dwc9uPIPTP9mhjovApwD2e/p6LhwFm7bbbKFPYN3EGrBlq+QOB5S74MQAfGk38Yxc
cA4oUMN1DubEFI4fUXjtTY/nPcYlP108oGa+ocV9zsnbAvk8gKJGAtrrbbSd3EN0LghwpnangWcs
MfqHbOK/Wc7bfX1HmPPHSY5RP2cCxzYCd/zTWTKL0F78Hx63RaHNRCMCyT+8ApcqyTV/9nfb7eMu
OP8FPg8rWyRVfXna0wab7qW1iXbZy/vbrJspSedjACnsg/sFdmvnB2E32eCCsPzjt7A11wN4Yf7G
b/j6SylqSiBe87Qh7EtFCU+tUZowciTSEqot3Nv7sZJiIqGK8xAa5W/L0Xca7I8GkVxLWaGpTvwd
Id5oegdmy/VfoKC18Zlu6XoYiYT9K4S7Og7xdwdHNFjXFCej3n0wPQdpsjkI+yWCCozlNV4Yt/ZQ
RcsVnH2fKxclh/OtMhPfkFs0nk0OSBkpO4ZydvhYp3ceggBw2CvAWBmksHx3cdr97PxZhJHWiEnc
gM5HdOKmqP9bzbBYyXPiYdvQb/oAEqEiClZlBRBdJSZmHO1FfaIDI93Ub8hqj3HYUqEhCDUzPfk0
Vp6Jg5bnhVOiQUWV67qkushbillhnmoVxFTy6Fii4rUmpUxgPf5UalwgFzK7Sd7qx67CvFc7i5oP
xYTg8BXPaswNgcG7kaBt/lNH4mF+d6HQoAI4MiuLwZANPlmudEQ5V4JISKGXaDBgIN4dsOhLjU2D
uT6XqjzX/GyrqmK3wSBEEeQ91ZUOBBRIMaRkvKHO7mtwH4qvVlIqhv4yDJBQs8PbFXcEh22bXc3h
wIsussMT7YCsuaR/V1laW1rVFAEN8YJEW5KOtcUwugfuL0+tcYHExvZPjQyB31HG1t0wx3Mm3/N4
oiQp+gfmZd40miqPzycLlYlXOqL6I+7xlYd5mC7WGIkOOWRHizWjs6Qde5tfEyAdudIzBqdCLHXC
uoPcP4GjemF52yltrU0Ne6vXIW1TCxXaLm1cRecdiQJ+fw5KICFj8sMNKHQe6kgBZKA+SaRn8N5a
c6ObGcFbTAiEhlVqatTChNTuelfCi8oW3VKjs1Ey10Me7vSl2lLJLJZ8tyecoP+CtFtrXxEoFQ6X
hD0O1QrJ5v5GQYqAS/VUm37JNLQKR+qUDittxELwN/agZisiHH4NChnGapw5TJXprIS7WPR9KcC4
lX576GaXzaGHMFcDk1f0BlXi+iOv8D+rqzvm9UJTuhVEW3M3Au9lXLwH4b34uKD+zk/6+4P8es3F
fdI/zYCU+ojGHiFfE+2zba9qSiajomDlwSsXq7WPuAeFTeFY4VRLWlGPeUzWSpjojtX2M039tOhG
dZUAirGYoys0YStMIWIkFW/7ZqCC0pD+bENSCZs4gsQxNWn6OQwgJccp0ZFw4rnPexamrj+A6V7S
iHg2DZkZu8W+6U5yIMY6KpUuNiDnhgZQacWH6cVieZzG2pHeqwm/0wAkya0jvEHpJk/wHlmJe3Lk
3mUEwGq1BgH3TZMSDW0gsNk/0ecyAd3Apv3V1cWgQJodisApzqLHx7AZhAeMR5IM2WUA88kVj259
JMTWtLgjq1LuM/eWFWq4KKq5K/jN7y9itXKx66cMsEJycW0RbHAHmjdgyB+iGsmem2xjg3yDDRq7
qoWIGrowUMxVs6WqruNFkdrBHlnvesHBpgJeKd9NzGsXVu2TjJ3UiLZzTGzRMXzcA/DtKV7uj+cY
48at7qDOBONAmMP6olTOIt2LsPlslNYom6/jk0ZOrGQgcya73ODusssSCsUrTEFdVQRCvFFBvYKN
1ce8MbJb4yxsQBWPGEPLChxNBw2sdWz/Xjrve8jE0K1doiWwLtk32SjibsdU8sgfR7oSMz0uVQNT
k9hZ0Y47oDDjAhopdinJFmxdPNBJJGmGXhOe5F8kCJShK9dXejSBNesvo40ZVOZyxh7jafxvutxD
3VZpkGnDk41iEBEMJ31uyUT3JHwR8VEZx3O9UDjrZmltkSQbuttshNRVyLHzle3UQQMDRX4w95kT
vs5it6AyWiyt11JH1bQpXnDdF4B+uS7yC1xeFr/5MlBARuEkQaHiZdB2WLCrIgJY6kkxA8k3NqMR
cLBZ9kBQOCQIlI35nY8ldki3XOx8+9Zi6oRURKOvqsuEO3TJM9pDWQ1YzTRw5swjxJ9tHcIE3IY3
PN5C+8u5vdYmcR0aqDgJ6x39DKM9H9WPYbUTGNabKDOPLp2b4D3jGHkXt+BNmIyc/ImANmVgChrU
OLBCRRR4M5ByHyWSjIW3T+mcXlmxPF94kg4nUAojOPy7DDLXKzu4JYql3cMP3ii6/wvyrD/ZAQ+X
65ZceTbqrUKMMeCGWJWg1sGI6h9VH73lDeerI2cPGu411zzlsj5MZfXrhucBtquIumEX9UHzJjO5
iZgstia7V8vwe8AAxvhdg2lAAwA/pg88qVPfnUzAW9IPlO/nRHpByZzo/OYOCXPlqQOmKMdDTQym
VAtaO6eV4La6iHz6FLRMdS4csjSB0g1lw8C0s+tGWZLT/8M7FOz6OYAVyUuhNAGtd0NKEltmqg+/
noK1uIfUTTMWIM3IqzET1Va9agn2ZYpP4xOb482pXCCF2obfon1bkQpXx6w12n/0IsP3lsrAtxNp
kRqbIDumOaIvsgXreZ6htkmY+XA4N0IAVVbCEtebIG8t1l7eTU6MlSVC9JfMu9J/nuf2n0uld3xG
e4zcv0FJguMTKoGw8LZHgMaTJazA9OOjayQO/EYoKB36Hd9uRLfBBBHmoE8pzFYS75Yn7iBImUH8
nY2lvP2jN/dDboEugr7HsEZ/eFM0+/O7qjsGkkuxCm9J27NwDIdQ+1TwGW1fhUopC4uUZw/FA3Xl
qrQfZFiWFUP8n9V9fAPgKdQB4CEgIC+83VgSk4szXmLnroQi4iZN+jookuz0O3oMmpG9SlenK8FO
cd2xACcxvmGB9cj0ZOHshXgFmH2Iz01JBLF7muaAlL/U3XtMASu/Qg0UlXIU6CtEUpywkuM4ew6p
d7bOxEMW9IjJ5dFLiEYjFetlHuwJRC0FcAH8HtDL0ESOP76iPReyQGb6wWQ+1U/M8/7juPFSmixU
Ayph63bPmqml/GKwzsNfWlArvFQNmFFUSTXZDf51EN8QNDP35bfjbcfjuQ3JsIBqhmmik5uyrm77
PcFEAlZQv6bXLKiXXbdgTqlqg5f29SwdrJiFsfQsFS9mFg74wEfDqfnXPHoR4EFzRfU0oy7eefHM
35MUPOMtrHDO2gW2w2ZXdK4rWJJXz7aV3pXKpDVkdWiST30Yfddq5po1yf/PLZCBTFOHKr0/XwbD
laeBzgzJPKUCpI7JLUjM/fYgMIgaJXkXJrKApoZnwkpMhwlQjUoiue07dPiRfF7NV99PkqxYaduj
UXrTU7eul3OudTNPGkSNrNywL1K7tf0WDjlgoTpBLXYUnaXPUk1AhISUs3nyDgvVGIdE4RqiAbwd
+aMDbSoYg09HyJ7YeNBin5c0A7Xay2yUGYj+oksZBDEYFERJScjb+Mm5I+st2moFk/dJYV7ZI+56
H9EHYUVGLrGoeyPYnTTKuswgmhfPBfiYShfRMmWYcRDRFg1Pz+JAX3AuotlCqIR9wHna7AjcYeVp
V7XRHN4GwR22YslNiHAPXlZ73d3aco3mpei0sH6+GPHKLNmP3UAF910Ld2OjjTV9Dg/OBpA012yB
ljvjfpKeDTE8adZxxjX/0DnoRd0EvzzEdxl6Do9o5olBKMBS5rBVLbqbVfXaK5h7X1MJEHWXB8gw
DvTqQwGT7nVz3Y1ftvppnU+urDMkqaegBE0QiRddYLETIDJuPRxipjhfqUt+PZtHAUsJUJ+yZYwC
pvYKd8+4TkKcg72+VFPzprUDK32gIaO4C+PWnNB9+ObYKHS/KiD2w7OdsW8DtsMkwORqM+5ft4rh
IWYX22nq+Gjj+VlfUD5Kb6yZur+wM1/kCmlwRrx+sUKUwfHCmzAuz95MV5qfiZwEYhYgC7b5swbd
3RsrAXXXHuGFmF1YPuqhftGQ5w5/fXL44/gErbVC4SWDBhmG9c1LowCoaf/ZV5qDrJYWIW0jhVjg
PNxIjQCvFn7O265dHvsJOjT2gI+A+CVPUpqUUfS7KULg2o3ixmNFROSUXzfC+goyH1gy7Mh3T+QV
EG9GGV735adZCTTYTtKlSXy0k4JrpJRepmL7VubG65M94acq77vlbJ3AybvDoipVZ216siodIjKV
fVoTMPK7pROSmY89iXIw9uyhanum3UkQuGeWhZ8ixm0PF7MedfKia87H3vx3rFN/q6Cqm9l5sAxt
a0AIXtqaIsDcoil+XpP0uKLKkyEEu2XNrjo7/sJlxa9TlM/hU0OfZgBEgyXRpv9HB0VNSvpA0uE3
qOgiD7U76t1tiKhZWL+YNR9ndt86bzNMt5EAcg05PRt7a/aSffK7HNRul14yfqsA3tb2+Ua8vJ7J
zkQqumTCREnO1gry5Kcj64SPvgt4e6+0zuXW6xr07L1B0DLo82hAgCE52WQqK2iIuwdWgPVcbtBq
7toDoLETWym9NmEMA8NWMqM5WMBiQ2BZLEPK3R+SFJX8nun18EikHzWat4CZG4NSAhpbVdGhBh4V
AD2lNA4rgBa4EDL744bT+TQMQm3wJbUrWLDSVByicYB7SPVnZFm4btgJNlKzydfW4qGN6uyd5Pjn
h1hXZcrK78EPSuJgJ/6iv6WzjMI8obezwQQFnIlOpzXBsAbbjU8L0PEzPLq2ok6Hjzaw2rqZh/NV
FyGmKA+80/PQvzI+no8D22CtMegycuQMFw8z2ZXabOkSo5sy4NtIoLJ0ir9tmq2a6nsZj6W8t2n/
R/fO/zbLmSXeZQ9h6YbdsceB50unhDBp4AUeGTNsJTlWQAq025cKFBxzDAjYEI9h7P1RFVcG6uyk
LGPpHJdaZgWbv5VO2+QO95bC0FWtdGEXdz0BeK9IjOTYju7fQknyhXHlCHCzakN6cPEduhgk0him
jPkgleBT2h1Ek9eJKKOnF6TgXo3XnNR2so9hcSPJkBia0vYtqP6tHQpRyyj/6NoWKRdGQlo1YpKT
rYCM2zOVmVhptP6Azv2DRih94Tfns8LeqJ+PRLtMnwrlNV2Z1/1AHp5D2jsBWabn4bObjNoJwQU0
FqMdQvSYG0qb3Q7Hw8T7KeulclY3RWiRQ07EWv8FhsRzdNIQKe7bqYruI5+KSNSq8KKEF/tgT52Q
U/481Wci4htwYzAhEUO7wY2SHoIbamEIBtRsq0Ow1CMFU2ErF5LbJMPiAIzRWQqEe7QtChKnlBJY
S53ut/96W0EU9WLDaJ+g8jfsai41g8tDp/ZAPaXhXCDy+DuYFljB3Dm7CgO4iur/HJjpyXGZMRoz
eug2qXrYhcBeFAg7qwBcJsjVAFliUweiLm6IGM8hwmRT3Z/MgA4BKaw5uhAd18JYSur+FPPZOgnh
NrF3OVjN2w56OpKJBYTG0i/LMjHJNvO2Mm636KCfuygLh5/gUw7VWbOEsURbMfhMwTRJZkG1uTfy
mYi5A2ZnrkWp6ky9ImiJHWug8e4tkRG4GIJ8+6e3KgHmMvRP2PVTembmBmNz92KlqgLh8o9Guj59
Yxr6cJHSI1PwkiY/Ucd0QvYkWUbpeLHg1rCVlHzR5mVuk2XLPNlB1DxQMslYRlYGW+to6QliB+by
iePgwxhvd1Nk59Yl4XKG8iKwIIiKao6w9PrItWK2YpdF+doFwHMp4B0RewBySO/B0hVdTvgDnswn
o0bNHefenMUcsEG5bidBgBo8Bu19/3W2EiiemHpUKx9PNw0tdqbtl6FCPNVlhWv5TYxPajGEjrV2
7KpvHBQM8uM7WOS9Zv0RmbheTQnGF70cUB1wezIcFdT6k6E6VzdtSEOmpPXcLLzzOsZ9+0uZk9vc
HLrCdwnOGukZXnZNKrBSECPafz4Ca6c1ihO6jWeYuvrJDhxd6PAUfNCfE2p1O33r3egVVoshainS
hws4WugWi7rtZSyXtR6IicMhKInn0Fz5+IOEVNMVmLiH7hgbegHdtEbrMqYfMxD38Co/yF/wxVD4
2Srb63T1EkXeofmuNTRGL5QfJjTTdOnuZnJ5TOg3r+06rI/rbqgzD2jI6QgbqSC2oDGf3mRwF6Qf
1JpGi+f7a9e5vY/x3S6CqNCpKyEAhX9tLpdLIVxJQaBE5DS8aSmqUY/kYwfV0SnyckT+ayW1MMvE
FBbM/vgqflrUNWzfEsX6q5Ew4LBj09ZPptMoVUC2v5KpWFD5nCabuYlgKn7KtsIMNGq0aG2CQfl6
mLTbncImoA7D9MD0/Bu93k/5jBDV1A6YIrbpVXsIbt2b1AsJxX954bHvHidxGwp6ZpaC46KauLRn
Ebms2Clp3vRbPv7mXrqniY6Aw1Dga3aJ7J9zolPwi/CtEZ9NRKe1PMGLOzgsSlNwy09daWdeOBE5
B7wtdXp7PW2DCQlWC6aW5hYXAe92SJzqmAQZ7I679HVAIm790SnCLcjcFusmdrQFcX5kJ01m0Wll
3qo1zjoyjmCXTQwOgj90Z4VHB+pnh7x9A0xxoBgnKwg7N302hu18qoxrVE7IfmmLRxLu8t9zgYOq
n8Vk5rfQofqP4pRWDDhtCNP7CkMcR4Pgx7jxEuRkBpR0L+gWx6iFvx1mvR8VbvFmjkrh+mxjUods
xhBtoHPeM8qvH+SvJ1jUOZDaeszb+iNmWCILemGgX+sXfPrPUf/bw2ge5V3Ssrrrg65oASU/U165
Qe3y4ZcpJVXnJ8x7DmOWi1WYWmK0+wSmGS0vn8LSTxiGfwREBFEykzh38IwzTD3WmI2wF06r4z7L
FiTKVVSRJctcuBLJPHjk8l72yvhJu4Dct5ohiEFURq5GbQ3fgGe4hkpznzt77FI3v+sB1liB0XiX
R9AzU6OW5da8k9IRSI0g3fVWw6ZMlFOOzg47Daq9cF2hSpxRrfBaUEkbE3fx9djIY/DS0FmbbN3N
DwbvmQYRFbQ+Ux2k7Fsk0wyk61/0evYjXiqLbWis4J04rWMQjlka/RLrHU11NCMpOXsZIF9NGAB0
2JGSzH2vJRH722YML/W0WSHNg6Tm9da7VmuDacvLlsdt7isO5ZUzR41sbnWQS2s0ccnd/vp8QPXF
krBKXtgVQ+1jF3LDsRJ7y4kklEBPrDXnr1SdOBRe3mtxjSO5XomVVzPSD92Kbvjz8YFHYcEoohiY
oSDypKDzu8pbFJK0Kftni5o9ZQ/mMQl5lJG+6wtTpBTGHRLcVleI7bYBfNcpVxtQtq3DZfJ8mRHI
oZgKl0etT2/93Nu9fGZ37J/1dmAQnNE1UOD2QCPKOMmCAkdgYJDxOa3CTfAet5StC1v3pMS+51mS
ZyTqb+mi6j/+joHC7KQA5CmjXqRdbZIaIqDoEZd7voHaayyIhLInt+6NWNg2CEHfM1y3WUTR3PWV
eploNEwMY6Qqp0Xkzfj9lLQz8pultKKkR/Q1JkU/I3+cbv7J2daFYXAqZWKRpzkl/n/BFbhUBj9U
CdZz3BjcrpBgNjntzaqBZSe31eDf3ITjrYUNukIXlfiYRhUVVkC+8ERJuIiI23JivwdgmwVekg/d
pPLx2s2mskgIceU2do44YCUjgXLGTQZFjprO8tEArrIArNM8Exng41jXegAsph4zrulq1lQP/1uH
GqIXVK/bDshfigk83DphzsihylJjJ6a+EEQnACKTJwZydznxsDhXt5lxdz4VsQC/kH3+IJGFkAtc
kndQZfwY0yYf/EqZL/E/9FybtCjgGTHngu8sTIXhzVxKtM7a6oiyHTZlMp1rfW5ry0euwkMs8fdj
O7MpVoA5UWPoGvuY+MdaN/mtyDwSGv26zOmj9Y4Ly4kyrek2rFumwuAI8IcMqWUfhI8dRZtInhSX
CuAe9mhy/Y5Z3hzKgpGf7XailTNINszbL29P75olQX6YJvStLfjjwukpGPtCBUR3Jl6Vzm2gAz5n
LuY+enNsAEBC2HQI6Z8fRlJ0tKzXDp6nDQF8+IKSC0wXtr7BPkC7dOPpdMffDHKiV9f4ec+TMZyB
KepIhp5W+JUCDUBcJOoIckPoychBtxMQdSaqe9irhNCHzeBJMqE1hknm6ss44ll1xQ/JcZ4r/1VA
PDJIJ9ZymoGWR3Aj9UPQzrHSkBQgv1CbbXPOBtt1Bv6lgS2Xjra5wY435LOYLtLSrKsttqdY4z/d
nPcHoMre5n811jtu4WpJWKAHmq53G8MPLfwS+AFzXn68L4bV1PvLlfp5hoxBucUIgcU5HZAP73tn
E1xQRWAl1CaVwOOWFlHljlKMH7xfbT5HXS56TdwTR2JMbCAU/unuGDNNrow/7jGv99I4vB1hVKA8
Q8oUlEhOF9m+HXCAtDA/ChBdNgvRIF6StLXbCi11SNIpzr1sr1AK7FZQjLjAs1QLVHb0v/d4bRjr
935kSmvwC2WURm3jOIxenSvHw/qv4AMPK83lF/IYay5fvcRVEudcyjo4V9o06xFweNH6PdDaCCvT
oS+SFu44ml2CGkQi26d/nV55qHs9Fawzu0hgayd92A7UueBKbuwFUhg+iw8UICsXPZFvxcggMnLN
hzKE1zUIea/F3g4s1USG2VYcv5Wmjudi58vlxd7VMxBPVFOwXLFDO5Iy2+ixPkFHzGwgvS8kMhNb
fDy5f2Gzw6iv/JFoJgF96XVCKp68iQi2EToqVoMaUKjshqkljS32h/GiSyhyzIaWUmPmn432l7T7
7MAgakXvrK9nZBporVXtf+W/mWYFC7GV8tzoYBpn5sUn8JX2bsesVj1TkDA5x1Rc0Yrf70TEFHci
WTab/uzPPH/jBa40oc8YvLRm76PrjqPs9vweuqcpqDfzrv4AjPfWJxYSJTEpJQtiNZqItRZ9mAIg
JIhvPi9e0XrA67PokM1fUPF9Jyx6PAvnx2+bEcJM7dt0FTPp6dMhVhb2fsgtUcOADa9r43dL0s/l
o5zDfwhbkYTRerTmNwBhDMCetbTYpsWUIV3hyIPmj7zsBkzBV1kPdWlLfDJKCMjHd5Km1sEREq6L
i1MKXzwNn4Z2szDCmN+w1nBf8iaCDKQKLsqVpEEMjJ4xKuhhT4Jb1Hs1FAceVocPKKfTcxzd04wW
Pj4jmmju87rmGytRB11uXIrvNjjSAfYWquL2FnpPfJJBzPMAkWgHURJdU01JUNlK2ScPSL9M9Q8+
T53VZ0OafOW3woM76q7mBAKoKJn1iS4VLWDgnXk/G054Hw6QS5oy64UzerB8lCzJuXx4aquw/SmJ
8GrEC3zulLZ6NhU0hhSXy/VRVkF3P30SBVi948AHYjiYY7rcoNLsAk/TMT3f241e5b809p8qL6pp
YOEJwO3JFAMITLXhj60pQuI6O3HFg9m8jgcW48O+e9cDdi5QMLfNqW7sp/rZp6+ex6OZ69M9fzMR
glj/jeX+vHv1zWRMJrhuvWC7t4tXlAx5MAR7ajmUbrXs80YdzR4ya2+2r7t7TsWegWLo1SDUtXn7
eU86CbAyEHXedItnnDvCNKmIUMMtWxkVJN9GPx7V/Z4eP5OQu3/smR1bftbfaxNeX04RhgUjPG/Q
oNJRvYPmyvmNJRXb6nVMoC9455/yTO4CZvbfzWwQLvyemUoFmSa0MohWMqqe1kqynRrLpQSdvB+k
HtAo6H1jqQOUzxm7rAC+evlrLQM9+AeOANhv7Y2ctT9mxKIgxbsH1k0b/slYFaM5zU34Gef9HAF5
o3HJQNwJQEHAfVzUyQ1LauMz5bJShZ8IAXfA4I+/O801inGGZa0lnGgESAdvRDxZD5ln8DujJaTf
8fd07/ktkObas35BI3zZsKnVXQC8OUqF/qyYOIFDANi/vYnpRksDJKTdJY8V34DuOdYIY/sjXcYw
kvXZidZSiYli0ssybkepFzuwT7lcBwF2tEbrgZLV1L76mvOsSEV0Wg1WMLEPplD047maa7WxCNM3
wnhroWWR74HTPrG1joui3L3zkem2JYLYIaGVV2skuCFnoTx0nzTwAmkIkfdsoDZLnxN6ERne/UyQ
leWnudIEBeoVQqQGrRBKoYvMkDdtTa1J9mfxB9mc2aVSr9+813u9FLPJN/ulERU290INa3sdp+Aj
xUjro6SG/SjgfIzqMd6b4vX8qsSju982XzS645tC4WHlo3Th1eKLDogadcdwFoSLZx/yYcvMsr4f
shZVJoQ2bv3L72dWvB8+9E92b/1LgC4ZwKg578ZGBUlzWMR4xjPaPcozwoxHBfjCiAvxCla96JYS
RxccARJb9AkTI9/qIV3g8HwZjiGjRCYwk+0pefqkkLDQh6TBFxhRPn+Rh1fBVp3Dy2g/AIAGWglz
SU1e1PYbHfqP1Q1ISnNEnRwqt3AkLYlhlfWR266IlwwXOs/M87cX3YMpNpjHJ+K/7LvMmUE5/kEc
zpObv6sKR0U6ngIl57kj0T3s630LDJeh/jGUhwp0qS5kojTaSoUqH+73gT+d8JzKu3TJyR4WRicX
sLqyBhasYvdVMVhpyXZVwCVKYoXJzpMIesqSSHZia4nVDBaJa8ulv2pKq4phBvr0jsYUD6CYR/Q+
ve95ab/UBQr4JjklWw023uuk+F8Emlsb4aQjnbcFSlSOEki3ruiWgblCCMo19+MgD+7XMOQPhukS
Opd1Awv8v7q+a7EsD/N03XREn+CClKZTNXx122YtGqAZGhVN1OhYWeUt0fbPiJcmOuBY3aA9UQre
OW/30YcarGgOhB0PNSx0tdBKS8HIHwRcroSlJpscrHVFs6UIzgVKBqZbTtBNXhpiSPLysodgExjG
3t2FrBzWpcRxsrV52bZwQKQ1EOJB92Y0izLn7uFvpI0t5DU+0HAmxtz7iqskW45+UiUIcDwci8de
KbAMBL42u6grodLF7mEvtqP/+KUzm+A9fjMKhLx3UG1qN7NH7t5phpHyydfAgF1hMWsP8kFEmoRR
BJkQNGKy5gAN4eQbvOV6FxNx9t4AzXBOe5G+z+QECOxegGfRcmcIGK7micCqvaCyutvctnblDlOa
7CajaIhn9yT97U9Z16psW/RE+uFZ2aKh5g9F4lAUHcJXipIgPcXqYrf+wmmvtYw8gwtgzt0HD+jB
lf+fQNyR4rOKy+LWUlPSz8ZOYl0B0gexd3K4wXDfqAnOe1+Zn0jyhYZWCqJUi/q/0UJgLIx5t8Ag
iXhoJvsNXN657XSYE2COGW3CXF0xzi3pyJM8HhvRCR1dq7nztIrOyaGo/mh/QDZ+XNYg58FDWYEB
x+5mwJqt7+zgpTIrc0q6r9J6KCmj7tNhkZcb0RVFei78wYOwNyYUoxf53yY/QFM95yLwKwesxaSH
iRr38PPjYhgt1eo1l8zPhSiENTw5I/jRHY/0ddeI0z7iomzDc4m0CYoIxcL5V0i6kv5HlnWYNhoY
YCWw/HR3TSiqlsGo+y+BLOB/6fZwkmWsLd6IjWHmORPl1escphPE3BWoOZY+8kuc5TFj8HI22P7S
PWNA/eGllup7biS99OpGgMHg6FDOeg4Ov2cSxSS7PQ83ggvd6p5oX0G88hce7MlUXaIom9IoEt1f
hUrbimc9h2NmgYDRg4RAcJMJcEJJQlWqUyzU8QV7N6C1GOFq0OuDfkTe38pHDZqrF/Pc3FKfeqoP
Uxf4lEoAwAs1M4lrkZca07Hbi1CxgOamOlw3fRXaS9Tud0k1y08o3TOVZejW86rfaR7zDhPGeR0Y
kTdztH7W3ST5tI/3wbHg8EdUc59IJrHg2xXzqdhhfSHb/iMmjLGLzunmsBanxSFTzFaZ/bRhFKAC
3dS4zTEPS08AGgX6x/RfvaV5zimqzX4O9VPzM3ZJWk07CkA4ZAlLLh0R63+AYx06nptz2pAj57gE
AnL3XliNb8TRHd+LvQRvPuNFCIJZKqJAuiP1t8DDX5f7S/zDTeABxPhW2esuUej4LVtyIyBYGNdD
GFgFk3VS4M6HPdhQJZ9t+OvlQRvYZ1EEI7DE8Gat9t96s4lBAzqcStUnvQUluatNbFzupxTXNmpf
6pmeUM1W05OZvlLi33Z8Uke7+99SVssUJR3BduULi2eb7mU+yFcbTg/ILUCoMAWL23Iemu8+84kH
s2dXQWgA4Z808Qs+ZFKvou94ZRf2X9Ay4gjG5YFI/ns3djg2lb5XD5g+UcuJM8rDeb6wrVTbwnwK
7xm/xXXD9v4McRBmCJRSAsrXR0f+xfoeeZaHHFGo1D2yXyhbiKGiU/cJgqOhaWumQOvsZYTTmpCO
9unXCIkZl820RE2yaTzB27sroj/E79QkGhL7qro3G8y/DDN/dzK6uuN5JaGmU1uU+WC00GAJtrXT
+7/GSb0zcqos/bTPnfNFNHD9bIheICSJ/cUpydjZx04qNkZW/faAOEO4wTqUsslUjqrPtzmukOk1
GyAOjhhc3a4STDDMly75Awu0O7gWaQfjdmvHLfJMp7MtrOc0R02SfClQrkni5PKIz7eKYJKOuFlJ
iqRGJjGOWAzhGe0DM51xM3wZYJF1B/3xcuVLvWqThtev28DhMPR948zweJyOxHCPWbswxAafGKFm
0M/KFc1eM1FYOSF3+mhPazmZTa1nSUeaVi7ZrRSpS146dZphRFICAZ/NhzYy01qJLQwdSCVbr9tk
/YNT44xFPzw7gCzBFtnLaVYtp6g4mquroihLv5VX7JR1Fc7+N+5zrAOM0Fk2Et0OXQWqeCI73+bo
+P10I01sq0UoSvkqZwqjz3co5Ko3JeuJnhBJJzprZpMC2c0O9W79VIzipZWFttqKeN4oQNxRghdQ
WeyOIMDtbDJPg7CVFWlmq+bawnrSy9ROiAVF49JMLVUXohyQalY9EHl1McogBZT2PtVmXGZHQo2f
VCcpOSbT+dftMljxajGA4+W5Beyi34YNrFKBSIs/Y8o3RLHwmu+FD6oauUTzMDzs7xjZnikIj+Sd
CrNhlBZZd3z+ZeG0M6uOGib2QR3w9oZ+kjKIJ6eFCkw9lt19hI+1EvW7daY9JgThNu+qvyciImY/
qF326E2d8jUsCIuIJTbn8NghMGzhXQU0/xpifCUqWOj2fZjL0zguJYUImrU6mLCT6IiLw7JCnvn7
enqelr6XavjHE1PIeKJLa3z+SDVlgXMPhKwt1u7vs9D6GeZnuth2ranUj+XsznznYa1gEED5NAXS
BVQ4xA1k6rWM8n3J0XL7hrtY+3RYG7wO4VDcoQNwKYCt+3tE076gaEMgvsHHL67XA3lc8vlwTxPG
79k8bEw2htm4yky2K55qRQb2zy47VM6eZqLF3hznwvvL8uGn+mRkK6TmBUKgey7ShnNJXTPkotPu
jJ53FNwTE4/QXwFJ34zV6TYw/4fqnOUiy8lPmbG8ZOEiHSE+4nFiR9mCR3QwFCDTp2RecUo0i5xP
B34mioMkcLyfxqmdnKwj/21vl32w5+s3rRNcq9tE0QdjWZtTmtmcre6rcSuYrjM34fwcbPcbkPrz
n/FDgggVfzhi8vf3B4J6l9x6Dy8bfo/p/bgSoJHCwq9GIIeyY9ZQMfEIdFUV93SkjnjqbEpv2elX
6GHpErbNmO6MoF04p7AmPnYUlAW9wQWyyi6pGshF89/qGetho1ppqh/eMPgg5MObHfHw+7pIaZby
hGOSi+9e8StCLVJC3vsxEYrDV+vers6qlfj0I4m61cqk4Vz0iG86h4laKaGVEO6KmqcG9qa/Gwpt
MZGU0I4X3dxeKlcwCqeHRDoEIJOa2dbaTRbS/QTVahSwWPOMpFFAiMj7E/wBKHZVKT5ieAhneegt
aFOKvzkFEJj2AtBeRP/Nkbr+y+1yzZ7dqH6lyPlasyFN9nXgNHkTe35mUsyTrghNTL6ZtXkBTT3B
BZpKi9eo1Bz/cf0ggdlkGtUiNnvmoT0Cj1nQ1UrvBYo49xzzrn7jd5sBrj4NAQMCJBF9BkIhOKJj
vqx3EkQh2qWpyDYjUYYf5UMLEdQTzcxyyuRmtu/THb2bT+sKWtC3Cf/8Dzpm4y32dZ2Y5VN5n8jy
eMnBzLWtjPAD98fLwVTvPiLJAukEoSRquMaQdAuEDPHeKdZciFOSHeNt0ahtJzlkcvmceqHjiJgb
SlnmLGQNDQZsEC3NhS2qESRO9b2NkaKTrF5L1ux7QSZcDjpH9tnQ62WTu7myOMpBnukf1TIeglEb
mTp60ZD+lBI00t9q67PSNKEV0feNRJIU0pV8etZd0arxB71Yif+zSAe7F7LQJQUNZ5anIje/RjJ7
Bknjv3QXJt4j3EUBCqmj0GEm4Sa9+n0kOOggS+xQPPwQ6rG6CUvScubr8B9ECObzK2ey2vx5rdhH
pSchT7peR3O2GBcK75kNXJnoFDd1ZW96IpXSkjYAj++PqO0Ce7avkHLJZ5eU4uen6i5TiKqJ4oxJ
VCpRNyINGCv5oa6R4nTfxpnli0+I4gN54LtiYgu3liEjhCUM1Tcm+Re3LXojEXPKTIlYkvUGDtF/
vT5V2Owse8juCFwjOaDDWkKAzhWTqX5I3w4oN55x5yK1azn7OZw5qtMp4h5zDc6wgegx6IrYwAV4
aH42WV3ch2Pk7ytKh/oRxMAvPQdcG0SN7ALUbhorLRPkGsMskk8YcyZL57tGbnq7eiZ6QXHJ2Jrq
djoeyG3ovK42r3doioigYHbRCNi5mV8Dk9zCOHaqcEncHJTWQCwDbhv9vU4NPx3LVUVdVZ2M30dH
TFdWA+wuqK/myXEjxuzMXk54PUXP4Xkw6x6/nQD6/89/wlEP1sRVunwvB5er6UBEpeFhzKs1W+Ms
QxlbtrL1by0JJDgw4jrKLKf90TFMUt22D08/t0Vajj7UuB3vbEsPGoPr03nuOiKvAx3igdz9m2mj
ybQx9FfXDoED8pCZXkES3QCVm2P5w6coEYQpyMu1NCpMVkbn0vd77Gy8k8z/jXvzNk7O23UNvSNa
TaDCNMpmAyvFRhbOx4XyD2nCqAP8MIPaSKFNKArJfgdLoDADGFytc6eAmmhz2pfsgeD7JKk5tHoe
bLwBpw7T5o/zqhLdV3C0WFybUJDSsMrsbsetWU5fZ2itdTlpyp3uc0L+KsWSbwvx26xDgdcwiIu1
YOS5i1Wn2IImz8dtZfVYYZS/t5bxq7Sck2BKtwl0DqZs0Q9qy2UhnpoXkSIMyERv4r81OMjNLNgy
PZ7s/2jjqiNtRI274BgqUYXhgntW0yVrMEmR6m2jfGDgqj1kMJmj/PGKYVasaqJZNxTVu0h25dto
bIyK5r016E/w4n2M9tKfvnV6BaVMTNTii1W/j5OZ9pOFMq2hcuvfi95X+uuZkrzlIazexU9Jjxrc
W7JpD3V6BQp+8ElbVAOCMglMXhKFdBGHJFDLSHaZx0OO4RcIcHYDt/60I/ttaADE7b7RrDbDPDpe
IaB4nTKsSCtTQnpM/Ob0kNdS/d3s02STYMo35pMeJyPZIWRds7pGtGpzHD10VMu2xPex53lkt34z
DQtf50fQS9Lb/mziDdCdOVBF03mgnxqUkJ/d19E+oJ5M7iYvjrB5HIcDsWMIXPCLKMYBUMr57uit
8fhrM2hU47msOjImcMFdg+05zDTLJPlXFOubnvM1D06fs25BKzG5PHi2KrBUS/wZdeA4tUsHe9QV
LFk7RtdHdiGnGNv3vn+sXGUIeoT8kW+0/vpFZKPxoBmAMDPV4butF473AL+U0fgbBK3+8TonFi76
tG7yUL9NHuzPgIUZd/oqqAmRsWDxerTs74Joy6l0jOytt+Cp234YD5ZCYf2cxz2O7Ndg93LqnuI/
EJIhCjppEeHECxnBC1THlbeIT2XQXi0X9ogroWMaCkHWs5BeSxONn/TDvkb66hPKBSjTX4bFPPnK
zQgtvyTKrJuecXin9KOnUrQiNBVLX+K9Fqy5ay8YJcaDLI36zCbUu39FQnrIHs/b9EivnPUU7lT9
YL2ohAR+Ypc6aUM0ZtMPUjWMSgKp9icfphyfplGocX3ayk5eK+LSs8M5+efCwjhjj7e4uv4kHVpE
H0ze7FnFi8161tExS/8QJ6PETo64xG+D+mhRIJ92BovHO25N+89SkSQ/R8Z6ttXidp38JoWXVUj2
DAriSNoAd0EQW9NfTiMbFPnirYH2ok8uhCJrifYkcOBlBvzp30TT1xDWpSS5XQJb7vVIbbDHppa8
Pmtv102HRoOfzweeIETJBdfp6zYsdE2sMHnabngTN5djJYcA/yMk/OGo4XfUxSgWH5/hP2i4UeqP
ec1t8V9/tz+hGlUyxNzRXRPbHZYXLFdbAvUSsE8WjX4Ceq7kNGlO2hQhnxFn8MAKdDD/pl2ESR4V
NDxRZSDiv9gORi5IWFzncQAjvqCrVlbMKDrsfLRBRkIbiqrKT3TTjp8rG9UKfD8L6eN+ScUGhg0A
eYm+d6dIJwf2LuR4O5XsoPV/O9B7pc5LoC+cqbOuLiiWRpAvw3Kvhd1NokwUSGpTzB/27v4/OpNP
pDKFyUh9x+AI7vn/JWOwg/6xpq/PJ23eaOyL8w4/TQqlJux1Z7NfCoRWYYMAMoATdmH86dych/KT
XezX814bk8nOZqD5jAAVws6+MroRx1xFNJiar9liwtOJMB6vMUtn5Ii+GCeNTRn8SxyecCQGoav/
lxoc6fm0fnmxcPa9Eap6QhFN3MCxwaaZAD05iH0EDtBZmNMcy/zdDXNm6BRkaKOMHBh5F8+Xo5NW
fplY3xLaXj9LHkoTg7cuw9gNn5IdgLjfEtTVZz4EtttczGYCKaMRZhsDHSNPgFmDxA9UhSANjhFr
kXEIfm+EerSo+c23ymbJIAiv/hdR9ZNHlHhX3gNAlqvCDmLJX3skeS9dw8aR9ggwWeTeaKL5oqqy
/nzOqxXIV1EqW3Rn9xw9d3cVa3cmcPrW5FpA982HdFhF8JmiQMp3YpngJ3cHkPFcsUMCgmy3moL2
vd9l/mDDZVgyC1QPWbbnVfrbkfOQ9thuGy0VmuHJb9o4mpK2wGPfmxa5yaYACzzwEc7ImBNswsD4
fuuivtqjtmwR2kcBDcL/2RGNqaOG+uy+ra2BXJ8MAstl4xxFd6pCAyNNPAwb/mzt5+wxHsltHxGo
mSKlZJf7xvK4qJp2xz5wm2S4L65kyX7L6B/nWdlpbwpvJGcewjWu141IrVdTZTFSoPwOaW2dhp6k
U7YBF77pCeTh4TYR6ZB0KvTlvqmly0pP9lijx8bLqfGKFhwxS5HFdFD861elNNBq19ULWohno5zU
EEhmuujB3/pf0Qlj4q3EY6OxEogpgCN9V7Wu9wVYi8K8auMM04/TusiMioMq4CgQB1nd70MwEYzo
mJ3HNrTCOfcZDsfqjUneXE/2+HpFDLEZr5gkfTbFFTasZv0hPvktquRhH82l+BqyR5DVag03EWAh
gpA2XsU/xtPjr4PEOHxmQZX1b4Ufq9mjuR5E3AR48hHKwlVDdYzGkuSgvDX77+ezN6tAISBZ1L/f
JwzrQY18+eSOt9ed3JRQHqrYTlP0odT1/P2o48YjTN2gbUU9eAXYY4vGvC+utkIlcWcbbcv+rPvz
ThLdd6zDzgOuzpnwc6ciVG7XoQb2PQ5UvtTi9/c9iuICG4RTqnP0g5ZARGT/zkfhX1impozekI6K
zmazmzrySvsu6cpaboB3QWfHz0aXpUKP3WsOs3ftKbfn3UQwkMMQhy2nLTfhaodgUWfU46l7ZQTT
HKRkREEdXNafI1tC+6leoFBIubrzFrdJMAzZmW3gbLuaTbn+Li83/lesGwWHNAj7n/mVeRJNd6Fy
Mbj66PtLtudEJjf27ODN7jtn6MBSU1oSP9TLH19rMWRdoN4CtGch/jDbfABH3Vo6qcY/DvvOV79w
FLlBFLMY5dG8FIPIZK9+rNv5JOGWEDaJiWhVrcBt0G/9TytRk4+9+LeEb5WLi6MYGvnr2MifLuQd
FMwB/zKDW3PfSVbjMaFySxos5V2Ex2NiHPa/VjcHarN1F1gN7iPY1wVoDYa1pgShYFaDJxSUVBzF
s2iRW1kTrvGEjqhIaBr5rpT/Q7Oiy2s8eSxj2sjY/Usow/S4fWyG/dhpG3VraCAiBfUKqOXKV7dY
Usws46/KEML/4drldGITjXKAjvozlJK54ZnR4VZRdgzG5Of9C1jm9G+Cs6nu2t7w8/l7u1AXtyvI
LUa17+kC7/CwkcBjBqSgod7ulsI4iePxh3T5GK+FUlerdDM+otWnWiWYmsrdKr9O99e2DVjUcH0d
4fSRdGNCFQmq9IHtaXolcSotPSEWxzkezGfxmnFWHwInQDXCN2AHeJ/HXZZUtLRcgcSWcnu4LS3J
roGlW9szGTtqTE2bvdUvHueMVSSRCRT1wFgAOYrOIO1oaA8S/GV7WiITw0vnPo70XmvP6zAsVyui
GigPG9I07EPmPB3TPPOOgLW/Q8ZGiNH3OISAVSn6l3ESVLJeaSy1MAypA6PUfEmRMUjjkjPQa04M
j/DS7/h8qhDVA3GWdY8F/oZ1YdI9KExmaXJ9fmNemiW1T6DfYOATi32W540FVwtjEHhEHC1rK+Td
9yYJKpyu9d6ykeTRRyxrAe5oYWcDAyAlsUcg3PUAcWFki2RsjWhEnXeUJs2FOjS9FalSUsQtz4gH
Bw9pNWFHd+4DXutam9mN9imbVHipLEiFQe7l8v8rOQI73R6FtAfmDBPg/7U3SUPschrCb4KWiRPR
UKOUJWftKTadYPEqsfG9mm8zl9PFYXptUIQv28R61HevohnqL3RQ5jdL62QTmfDjFAAOOuaUEia8
l449mIb0RSyms13qVdJ+98xc/WKkcRK+BCa43FTgLeuLGf7SkEGOWUBtXBswFUXKpAPRCLLAgnX4
Eei7fdGn6n7NB4jmcl3f/TmSuRJNHwffhHDfBHbFp6ezSyWD9U9wlz1z+7ccJBT1nhc64+5Gh9mO
xN0zrOhBMk+d1wFm32kbvjRrzAnb28R0HV9wP9Scj0cLqQjHF7CWpE48ReeaL0SknY+5WwS91Hx3
FoXM5JcuHgzxS8qj13cUP/nC7py8My5tmp+cTM5VN36w0YH1jFbqdNGMvYqZPttAKHIJI7nyLx7t
Swq8cqcDLrpBMHw+Gy99Klm7ECSS6xPZdGhrJASTFOyhZXKZn9GdvZ+AJBOSVFNnlj+uH1pa24y+
qWFmfVtN6+KBbuv8vmev5zxAJTo5aZp2/XCNWD5IPV30unZWHwYe6eeyHudRXm375RyPv7FHxsFp
yEsI4nVxVTF9cIKrulTuBktZmgc4AdQKLgBZx0x6akvIxS4L88L1JDQaJP0PC1jliSrJD3k1GmFY
zSsiKgQn17J32I6Tw3R5VO/fd4jncWx9GuXeVDWAnTqztmEUXLVH8K8hG3wlculOmMGBMtBd52bs
+AE3AGIn2kb4UfPLOlOv2t7hn4oHGR9PxiUH5ejrjMu8X0BVKL/hd/H0LdyS3lcOeblqo92+Tsew
/sYmwdUOwenWttAyjLkUtG07rkS+AR7XW4uk466e5hPsLMkLCJ9Z3Vn+SzuaYikfNUN3fjmPB0qi
naFS9s8LcD9ZjkX03rgelm9ekzC4g7DAx2kndhlli17ba9BXE7lOMYdK1TkuVYK60lVkKqt6f1CS
W056rLuOalfGPAj85EIEPT5GJpUvrecyy+uMO2z1CktHu0PsqNAOJe8t7npsSqCp5vRz+h/kdzvF
0Yb3XVm8wfHPnwGb+7ePLJ0ugpl0NcxI1KEKLAc2JH3z/oL7HtsCqWLblyd0Q5Iw6wZ0tXJ9MGV2
S1LddXSiKzbg2co4LW2ki1AIecPDC8reNT+ajt03LwaEo0qOcdLqOST/Z2DWGGpANoiHNjTjM2sO
fX0AV31PQz05sUQIugy5x+FWDIDFAFpwmzqij4q9xObBd4xDX1CpKiN89PVnKt6K0akh0UJDpvCB
EEn/dc148p1fuCZlWmxCoy39JyglGeu5BeAAcIRpy1PIcn9l0HmEph+4/WuZSnhUI7RWlpt+Vy7o
hFPqsY0ETVwiu71Zkw+9Ok4w7QlO02vHuICzRsxDy7AGf1o0lxH8Rb/G1jZT1+lOeLKpC5D5svHh
8uX9ayYmrnpOUmbb2xRrxNauobpKG9NHTnG0b7BDfkQIay3eWIovezyph99F/7j+RymPjVjB4YMT
UIpThZGD5v4HX031cZWHD4FrNje2CB3qSEVcu/yIBgUt4ZBMWq/IXCciMJ6MBrLgh4pr/MlejeXH
stLJX4kO5wcv+JQoP8EDheJCDCR96/V4q+LX4080RYXDcyUevMSdB6Gaonl0+sWq2UNUAIaor2Rz
QPIBzM0pQZ408aJ7lMgRLnsyuH7Lx4cffkAHPRTmdsypV7mVIcdjSN6RS2JOhzJluWMfJimCBFPe
WSMybON6Th1if1pQS+pxsP0nsWk4JapjEKH5SpRGqdCd7Flupy4tAJg+CzgrmV6lN21I9nsskNfs
hQF7kKyM9GJNGfh+o7DrZCLhfI83sCs8+L0JBvYOVurjXRWKRFiaCAr8nOlmHCcUgJb87A1jnHXf
uXwVIJ2vlVGd5zi9YEvoTABn5+IZECmKjGkin/wgXgzgynl75J55kqXqjN2R6+p6109/vinsXkrL
l+jOLKtt2dF13O8KEnuTCExMEmmMDq+eD/ERWJlRzWybdxa+JjvlQGFfHLGuJqytfSqLZlGrre9e
GfkOrApiUOds+nbdOGnEi0JOmQGIeXMEFFQN8t/XpwobeaPoqCEwD1A6BqI+P51mIROgrFRIu2n4
eIjcXi1fHEiotfmgCPe3Mc+ixi96UmM7KKU91OwTm0QTMyzvvuO1SWWHk0lDneVkrO8jMOEt1mz0
GyEJ+TZkNNygD4asPSaFiif9EXcpRAZuNQj9EyRNI/2ENVw8xXCPXiL2gljzbaYIAgMONUm3iik8
WCHA/rb60p+QhUYUFiji2mK33UlGmfyWz5irq2M6UTTxgNuePTWn+v2Y8RYIxgySZZg7rHws2LUK
FNbrdyvtzqnF8BRsxLf+UscqUmtd2SjfOtgDkhWdclpZghfIS13gVbVkaXbCZlEwyEGUjDeHcR6X
Pa6l4qFuLQj0HHWD6+RbOxs8QIv3PJoF/GcKpgkxsCLBngc/b0xkxLQQFINJYe6ToNp7mNrOcabP
YeEZyc1NPBsdooqJamrGGVlDdEzB2aSfsYGgfPPBcnPzW52WDrK2JUVlf0v6GhOt3TOre8zNGr2d
tDpVonGpQ7p4Y+InLTnJvCIMffqB11GRC9L3ERNOEMjyZGMyERm8JKsenFhmxFCpWlfqrvyuStx/
qd+Oma/tyY9oKiVrRo7VheU7pl4WocyZ8u87fAiCzz4gR2+cSo5aL1bqs1ejNO1Nm7W82LVtnZRy
Kv6RkKX37HVloKLeRHnF5FGiM0oIzaWFZZpCAAbkokvNO0YoFl/vGLr1HofaQEo2N1UBnYcgwQmy
dDeDe2T7knMOv/BjrkZxpBa+SyK6zOtMbVrqcVeB8NYXktu36R3OLupGdqxDzLqDPfnWz+12UqVP
R5AiTy5MnayifTKh/1jV94JcpAGgRcxyu9TVAIunUyCb68r93D+iAKgfw9cl8lrH7dcQV7+z30LX
r75kKVQa8gJaDmvlU82CGVsBVtGu5QCsbSjaW0acmcobHW4c/yi5JhxqNp+5VRXTNajyrvRc+JG7
E64oUlZKUcMTvAduHj4F89zmEQdsnlrmRy6/ZC2KTqXt43UQQR84GaFtqxPpswryFBS8h6H9Ozd9
rTtcvJOJqW6CHrvIO6mWhWLDwFjx5eyW3PtnUeJl0Q5fblLuLw4rkTkQ89IsU1DA/jnGv3Zi51/Z
j6YQXdKTOJeqDcXv/0jdhWP8uRrvneE36NH97n90sam7xj/4FFI00bnYR9raOLAtkd+iBOjcxzIj
AMR7tHRdEBGw78MflPnxlRLrJekPDsOHl7jKw/Kl/u59Z6tnJrIUeJsLNsUycjiqIuXCgwbk4kyc
y6tB2dyngq6rJBxd80U3dsOUWEvK0Sqg7K9RQgQA5SEuqmom1Ep1C0WiCoMV2bX0e5dQeIaoxSws
oVfFA/PVMOHoLF4XrYsizcrrJbtnYqn5qcIX9sYHDsONOvxVDBWM7XHwFUxaa29zWV1taspnvod6
/gKG6mA41tg551ydJ4oczSOyMIvQUcwpkTDmfN8bxNA7Ew6+gkQkuk3lzzGPT+B0EjkVk+LfR9zM
iPp6kcZYHsu4GDhwR0we6/+Y0qh8I3Q/gUQEHnDDnF/d4DMgmqXOYcNP9EAisd6wrojCwjmrjx4n
2rlCQSycg2Awoi9pc52bdoDPF5PlpSR1Cm7xjWC9br9+f/gnt+s9L8iUqDccJgLVf2ZDonhGSjeb
NVICRh2zZLAzY0E1KxAAgEND3unvtigWlY1iPaRQ8ViEGzEMEvamZlu7e4DbwT+cdsX5R/SvWO48
DfvRMYP1iIZXXaS64w5AkccOtNDxdo9Ala4rqTUdpmuCqJ21bsev/6sfoemPHLckDg976byhuKZG
GDNED+AJqShpuGICjNa59/5vReH62OFy8fbF3czdFU40iKA3H6vOIgl0N6dfi7xMUli79z1tx2Ie
ilREcd+d+gqwdTQ2TulxAr8uQrF7hjrNz5FpYmzC5E0v16h0xgF4piKTclmAlMiSkNdrmXLIpDCj
4V7rYCIuA8JdzEyGD70W0twX1P+L4uCyfgRFCcYLJ5V7OcZw7MjLZeSc79UqXNe7kZu36EfOogfR
Y+5dzVSgxlWnFTNahGxDZb1NwGu0kG7fB9aGraMCLqlJ0A8K/MEq8mzwYLsb+roS/iE7h9YSuMN9
n1Kl3iGhOYucJONDyUhokGk47JH6oDCEQlxNm/6NNzJtD8SgWk2P6HvGsTikGeNORsJ1BloFFVqR
smw5Oq6B92DOn3vpd2i3rSUOxcXm5h7TtcaMxy7xNWcyCe7LUHyfbmImrrje0TltolnO7GBjaxeQ
LlXtDOTD7kX7qWVLYvHHrhoTNDq9I1POx6NMuDfqQFo5kYvF0w2fXf6f/nz0KdTaf1K2n11PZ1Al
IxmsQpJrqLc/sK53DhvFx3KusMrDVNPfPSUE0O59dGpmWufe/8OgUN5rQ0kyHhVW3oZsk/4TgYbU
j3ns66FMhNmA2NPLwkUAbRdh6lpNR1OCs+hCxQi2T5RZRYUkwxTFBmnHtjKWt0j1v3b7HNyxLf32
Njd/7h6eF39pc/SR4zV8cKbwtuw5y3gV9zP6jNySD/IovpUixrkKw5sQWdjoK7RpVn+Zy3j+De3C
5XU+/rDdYqsEEY9MUkVjcjAoUkch8GAYV0pFCk2Qa0NiqKTC1UohxdtFVWG0Gwz2a50E42cmtpXl
E7TIl5n+7xk4WsYy7jLBHtCU2X8xcg2uaO+7vwIzT7WtJ14PSqknYA+ASsOGfXl39mb0w8uFjyK2
dguqXMKsV7F1ATZBGf0ecimPkOTGzj/26kflDhB4hIq87e2bsdXcrK2XD8Id2w88uaUSdFWXz/jm
COu39dky2WfSZkN4ScJToDqwc9GcwOeH9dtFAY516FKKh51TBXBI3ndzz6P1SG1+uepNaSwZmIF/
O9ckOVqAzZcHY3A3o6x2VhEEzYZqZy5//wMnAv3zE9RjID98tdtKRetSmaZ1kTbe5TURhqUi7w8+
lL5mjA7ObVRDwW1IGM2OCvE0Z8qTljjmPHmj/z31ID9gUrFIsSyESDoN475gpKdhA2VREzIriA6J
OQv0ZNHkf8a7JRTjtBB/rrFLAScO9AF+S6aCRIfc7PMX+LZKajfxWqkc7Yd7yxndx/P3BzFj/nTV
kly0m+qv1dcsCS3RNHBMSZVEzG2e5itOunYV3cswTrWr+koQjkHNEUDKrh86n8rRo+tPhsYoScrf
YqcURV3XHY0clds6v/32mL40ja/UHsltG9FRXpMJ4ZPidCBph3aXNfwD1Mr1Hlh8bRRoodStOCxD
DBh0QLhACumP8/eWeQ/CyCXWpgHjR2um5s6YN02yEEV0a16rpTYVFgHcBds5FqPd/FYy3xeriCgx
zsyxD079GIhVcPMxI7NZEJrDmrVxXtVUAQzHfb5zpJcEDAxhT7uZMUBgwImlUg0ZqEmQNfUzYDXl
EgK1PEJdS6R8xda+MSLY94fK49HyEalZhZwYKx8PxFn/lFxAtYdq78ZdCnFeGWn6+R+uOhBpkZpc
w1RcoD8Cr9cna/sURcs8QIiMhBFV4Y9AnedEbPRICqZDY7gAyNykYywaYSe+ObKhn/q7aOeGUzPc
IWzno0m0qJkFQnH+XetNRGRntJ0tnESgfSpf24vrRVmu1n6CZwEr3emXimBvk0nZUZNH0pZHfDE6
JwdcP8eEw4G5IEPOt+kAxUTuXoP5RNqC7MRk/ZLZS45sKxSGCcu8lnMFFrZB0uedPL0pAiyNFFRv
TTJ/EbbR2/dvy6nB3SwiVRWncUNU3NdGVrSpvefgIu6o2iElTFqXDzTGr16FNPi/H5WZqmoAycMc
CMwLc1AH9AMjzYagsNsicvw+Q3eCcS6f3o2f2E0vgGPwzpMgsD+tAzfgUBy9IovtnM4srbShRg+2
+WKWIS9G5Nz+QSHkpJHLdHwR90PtTPLVhrKC4mOUgdCmVq55FK0WRbHWE9Zt6u0bcSe4PxM9io59
tiBGM7TCGvoTrG1878D+lxVlqqmuTZ2yLZmI13dZUuXVvHbOqacO1u6+0iDpkYeUZsbLvj5W2MlV
W5lHfkc6KhYRLtTXTQ0FAfi7KuJazby/z6n9GtUyrxU+RdgOypjX/o2Ygstz0d02VODshQEkwJus
EoJnk25deb7Ho4OaKEg+xDuwrb/ptqaiGIgFpj9nixDH2CWyfaiK1uAGxt7VWnconRIqjPqholNP
0+VLlXoqWL2gdtNEKFizKHyNi3l/0RkMSdl+L1zUUSrVvHhWhArtGfxISXAvs6IXpv+OhCiYnOt/
2DHxjPfGcvOfvyU7hs4wYGMrgvItPJTToemvs9du2QtKHhsi+gxpm4rDX0/zUClgopFjOiyikmFo
Gl4nedqvX1PYwiuvJGE2Q9HMx1/5EiJ2vuhoPrJHpqD40t6oDD95S8qrtMvb+JCPxcURO7Xcqkba
NQLyGA4din6GyAO8wO0XqUP1OEy43UvcfbWetPX6MMzbzrtGJcZYnOT5gGbi/bwh5Oicbc3lI3yt
jQTKWo1X9GUNKwxb27HtJkp6lrSRU+FqL4IeuPD5xJAozjX+1S6GvXnB68/P34X1388vy/1Tk/7l
Jj6wG/MylBc5pxl7taWOPj2t7lv4+RNTHucmIvfaxrUkbM9DPtf2ZeTpEFhbJM6yfu5OmFRAgduj
nITNqROTds4aG+srSzN/NiMfQta1XCpCjDwsrToyVccz8T6wJFoJ7NvN4WZlr2ahYzm2RftAHRZQ
spY9msTVwpfcj2JwFSf8V2oF+rkIpkpVa8zqXN6BBAOmiNPQ1zYq0qbfmCCCMtK5KoQsjqYxCKvs
dXEaJg/LYY4yqKQ+My1/oKYIc2famVxfHtEyqdNXi5uXSLZQqMWoteMq0n/UxsDk+Wyh0Gu+qFKs
XXVSs9uF8FwYltx5UOoGWyAjJZ0ANkTmkpuOWlUM7ML7B7BqXJ9e0Lg6cwvgoHoXFwUBfT3tvgSI
JOXM9DJ4/6m14Z4sr/+qYgW/kktljffgjyRYjLuHSZvgFItAbZ7k0hog6W3VHs0gEXOLvgdqsa+T
/7zATSnZNARnbreMhpo5EV44YHlRZwdggVgp1nM6Rh2Gg8VNwuNKDNiWeapHQtoFY1wtvcl241wQ
yMzaEjAGIJVsK70WjRy6taIXcMvwdz2FFRJ5b3qokznm/RTdSOMHqTObZdACiKm798BdjkiMbxXB
PV5vMiW5HycvVjjqKAL/Nqd+h1u/DJEqOuB3MveN7Dgm06PlFBfF8N9wh6dPA3oUHerg/HWa38TQ
GWrNhYloiAR3dETuD/tVbIsGfu1zxP/xmLaVbJRwRHth4J2J6PcSTEb8aoicLlKqfbLDHb0D2wFc
M4XxYHkdHnsPWLKXJNTY2gWXyyPw2jDeVcEvY4hiLgWiykaUuon14GE8yQeesur3iG/oBOQPeWaP
nSg45sU3c0ixTg33v+/c4Zd7nStKxQsxrM3bHkZ6AszUuAnpA97Ev/5yF6LISs3XlY27BGcOGGQ7
uD6+OMwROQ6ySVV6UYqhkXBsePQ4vh7bPZ5A/I8Nsi+C6HBBuSJKfZ+YdCVHedG35Df3jrc+URJU
5OAbckLyZqPh+qW4CY7BY245zbR5ViWY6lFTsbN1ZHade6n7YphtTZFpJkJvcqnEigHljtxBuyuq
WXo4vGPkTUhkbJdVyZqvMedJp7cGIKThgnTNT5DBmz6wKqa5fPxa6AEvYHf9451Egxbhs9/6V69f
PBkEd/VgFFtIcz/dGsBCamKREcya5iy+nrQ/wioAmZpkgQd948ycY7fUcAI3k9OC7QfjzxSEY0V9
4EEIkiqDQRIgfHPGdFZtEBguXjR1Nf4PWpCrPGI3p8LpNhb105Vuy5iyW/fnmAuK3pIdWtfavnUK
XUZLf9hgnwavxsqOiWqk5yjwMOza7JuuGgbG7lTGGOLBU4VOwiw2sU4o6QILiyuRuiA1e3f07kWc
0kwqSJL5GYUO7BU4HI6dTVRwBfxtkW+3oYc/TlLE+PFso3iM/9iderE6QDyI2yixpnMypXQZTZwU
YYYcWrkp87HWF8++OKhUsluRVxBRqXX2+fW/vhQAbnLG6CIDdrKwHvwEamdctVc0oxHHtkDn6h/C
V8f6I2o4fPSKfpLCyycv07kYXpeQE6ha64aRNwJPjqr0/9/cQL53dwXUaBK6O8WN/AQxm6IWp6T/
j37C3lMrcgc/csosOXR0ILLZ+iXvEE6+mRgXdpOp5o2vlqUlvkPACMiI8GHD9KakK5yynw3wh+Gq
DYsp0NB/XDWkmdC1QgbYvVzsaEOLD4MrfkVniajFPwZFArxXjW4wsQqUfAfBWr2W0XYgIVHX6uaz
somB+Gt1u1diIS5rDrymmRUAcKvAeQgRFuyCKwdozKzSShYJ8Y2Hf0BTQL057k5ncweCVLgwERPS
UCsuP2J+FTdvA5HETZJQP32mKiUyj2po6hqmvP7VF5N6dqP3N000ttTCdApX4aGOH8wmBRa6MjjD
208ytXc3ptmPqIsXWfR8cOWYehQN3S6rFC3p0f1CO0Dq+lPialSLe+8zMVgqvMscVKhUZW82x94D
ebPW+SwPFCqE57i+FyZ2+7XqSVWbnMulldnBUkuyCIieciROAJVjkFGCxX48qa4shsPDIx6HL5fq
OZKyvqVDEoEgIwcSmOvVZ4AHW2X+k92q2tffTribFQK7ot3mXQk8034wNM/bThaTUKc06qYoBWwr
3MqvBH9QAednBwKDr8GQJm+yZ2cJY7+m+9eksBxU0u73s4sEUlGRJ27JV4+DE0acNiVFeNveC278
X+a7F+jjFAMVCgTgzdOk9nY3Bw+c2WtL5rMBueHgO6W/IjSaDSHAjci5ErqXWixR+2g1/8KL25wj
Xd8m8WmhFpMIjKPL5A0yRmdmcRZ2x04qJgcSq4sCCAifluQgmgMCzTnyi1i+geoaeW+aWfxyGrtx
2EcD/PxPDZ52gJBj/ypXnHoszOdjPIMXrp4xqbNQfJRD2DgQIsBBL6yKms20qwhYhP82Qb9fA62w
30AAN6ARyl2RByvtCqyK6otGBmevQC3oqfSp7mgtDu2Z9OVEBs5+/bau3KDrrvgFJNdK8WndN1+K
0rUnbfGFbWSUZYPfqD9/fVG3mNFabMIcn6Yfy8klmnbBNo1/S51zBqVVY5Gsne6qMOz85TsOiLeX
yoV5wZAWNQ9w2iSWXjIj1nounCysHgC1nqcSZApTLqfkY1w8HLaq0gxiL6DOxjryKCpb884VFWsl
Z+Q3O0DJJ8yeGXihMbrfNe1GVARpLHM00IaBtibQlAuAPx84LlTPlTv2xdQnsCvp3sH/pnFhTe/Y
Ie/S0GN+HcQxnaynwE9Pl5HdzLPq79teEYoHRwMnhshbqejt4nYO104Iy0EZF+neIV36ByNb+DHJ
ZOx7H77LLR1HnCD6p3NZhlASTeNwB1js0/Q0Pqb1aXpeosIlBVS+I3fLcQRCIgo0u/cI7h97jGyb
WlSFvkKMmZbWBsAOPnxMG0JxcH0OVAPqQEqIzY6Z13STIpm3Pbg8ssSFyXFC9w03+cYDovsuhlI+
alYPDpR2NFUGrBEVjHX4v+vgd/Awvwec3e3Ebu/Cgl9UfLZ0nOO6r4CNrBqRDl78Xyrmi+1zLkoJ
3e3UQDVDBg/PgdmAIJfeTlVw4xYCs2d4CzUfExEJKvJ8+riDq3GqYzpYjUWRo5yEzeeoSP9rHzJX
47e7W6KVMmxEmGahIZx9m9QJnjQAEVXOCP0rkSkhdTs0gYJuX9FJ6Ne992LClaDnD9q7IXHPh9Y6
mCOLThFxschHvB60w07P6Bm2B1K9RXB2qyilZa0ZV9swt8Ngkb6IpyHZAtCKVeYl0pX3HwaFM8C+
v693Dj82IoeKJ3q7LWyIGPDwnw0TxJW183siKQWNe/amPsxIS3k9Uh5NsCH6nE5rsf/VOy18Vlqz
gT0+q/stCdNm6+w1V5tMtqc+ypTKGyEsyAUMW7PeI76ilivJXuOM1avzIPuBq5wW4yr6dPc8KHQq
WHshNOv5BCqNekqxb0Tw6cGMgnTvITJvqrzXVzVUcyN3WkxeG1ww5UH2IufVgT5Qq18c2kw7ixUo
eOXN/b07ArtnpVJTTwUQqnroRsqCc3L8L848BpGyLoNXEBXvGHLFLapXMlYknI9OJ/UmycFQIU6p
4N9X84q3NG/7UCEC1EU0X0fd8MQqskpm5r22Kdlj9PfjCOqyIDlOlBPYCgvs+ANT6neDaJxRJG5p
+XNPK5xYb7pTKmyNLhJYAAWhTr0kJWJcnt9X2K+7owxwLWMpZ+HWRsQsS5aXeRcaFd0sYh1W+Xmr
u7pvR8JU9GlXvlfAUrzFtv0V0f++XKXWoYpPKd3QMRx/ljVYRr8C2E2o5itn8jU90V+iTEJtIzTG
e6zvQ2v6wP70wEc8iaKHYyneZnqG4W4UKvdKydkA8I+sZg3iouDG3NQtaHWtGbSmi/Ut/tmflXhp
H9PjnpD8xLVIvM3USC5mi50jJy6vCoJ1cjMsHWBjFblLwGdnh0+Uc7Y0KO8NiENv572RQCbJKTrn
b3R9gwH1qxDjZQ1MHi6IJH/51xOfq1okXno3pKktkVdP0r+aSi92ELmT7XR/L2DSa33m7vHLRTf7
m9ChuY3P6rkl+2w+eZ6RrSfvKNL589u+sdmJmGSIvcTw1cYM4YRgQw4FQmzYbjJXe5yhbQhqLXlm
PrxiIxjsu/Yag89GqU+0blfTSoqEtbqjhhzerYxxjHdy9TIbKd6hIswLv12n8tFVz7g4sNIcaR3l
NGkkh1GE7iEskwnXXJht0GT3MKP/nkd91LaDfQNwQFqICHBN0o2sVeB79Hap5vGP4nLnvfHDGsR7
W6qO1oQQlMd3R1J9t2O6ZKMNwHkrg7acxOvqaAHDlW3UfGZ8TxT1SI5GMX08dTxm9A/i3DSH99gE
66Q8qX6SiJasZ0lz+igGPz6N8A1QQy0n3F/YgTnpCK33y98AL3beQpAUH91CHUH3kVAFM3t6imBG
t29KlSLLdtnbO0cwgyUktMpKA/FFMqno7L7IprCKqKbBCG4ZAHTLJ0dz6nwi2+yFK7U/1j2+Es4n
CeTcOOUPStSjnFKoaCLGr4BMjk3ItZakcnScIQgFaHnJeeUNlHF3w1H1u0Z8jQFUn9iALyG40377
tL4cqLaoH7zZCPENudjLJsKrTn4Jb9LgxA4hC/7vCJCYJleBlMsW0nVv1tQpIElD7GVN21PUNDMF
/nfIy1zX8fDoPI8qvXfr/B4jq7lUu2u8wtt/8EFI99L+lVMSyLaqxD6Nd65OsnV17WEzLNQFdBVd
agIGpJSsYaMlucvE9Wf/JI8blG79kSMtmgY23JSNG8ZeSrZY6aWtu4dSe+N7o1H4lVfn6/L2VHmw
rVlzcyTV3sFcihoDU1Xn8pl5qeEq5yUtd78RF7aD6wFZYt4vdy2ePk/EyDhkmJz7ZQ9ZoaWSm+qT
dvNVWou2nJAuvZJEMG6eRmfHbuLUe5GmgG13rMwh+/dJzjJ8GGgZ05qio0tSBm6uyaAS/NeeXEJT
Z5mt+QnDGWWFS+/AhOy+ypvjWy9H7rVDgB+fB/QSSnoK+lQgtJxFoI4ZVPn4H9Q3lM+4csPNxcCO
iUKSGKEPqNQWU/pV7Zi0v/N5TXb8mjKeDO9zJBEY3ewrRPa0Mh0vfFiRnOHDAlz5qe2I7yM1urhF
cpvutHFl99UEDAYObc4QZrpso6jJojiENwY5xadvRLBBKdM2ajHIEnHAYIy1D/mcM+mgPIWxKDYY
2vyICOyhkC1nh5uZLOhljyY/xcJKaXzqXqsGoG5DTQRodxu6jRmoxSgpgCl+R+3oIjze9oJ7n8I+
oiR9pRsxq7uAr29Vm41ipd9jJUqVoOJ3khjQdR6DWDJgY+9efHumYWbzOya3dhfY2BV7ZIYlouap
VDJWFSAvMCyi8gNqYw6oe385/Va/qKrndEzZIcYhOdRjUsy1Als1vn//lGmKulf9fAov80KszY4T
eGiRmiw4hoeQImhSo9ea0NSFPr1/WG6Y7Hq+iyhw8MU6OsSOJaLdkYqhL5mpZb3k9Aw63Yt0aLGU
CFcELSNQ+0jfH6mei1NxnUHvpT3EYFgK0bZV9jIMWuHbmcTSc9L72Dll75t0KzRAEqz9UfVL0o7b
/tYNpBXzS4ULAIWkjp55CL4bZU2Rjf3yAV8ZHXS27EfOVpNDGvlY/T78ylMSwBGglsJXY+tDMrHI
9E2LiuYABE+mSNqyLhM2VkUiZRQSOglZbfOIyq9C++bPRGb17/CSumporNvfHixO7tZsxekzoHdT
DzxoC/TdQjv1fi2v3ssbZd2/vok95JIcLHh0DDbx81STKuITTBZSZHBWIpJA3rTIgCaYJyfw0hXR
f9MXtLAGLFSaTQeZxQLmDRn7/lS5wgFsTEyW7IHS+gsp3aPMsRmjIHJsSZaT6r8ySOTZUJsjDLSw
2eCabbfdqRpD1iRuWq0kKQoHwyGZvTtEzbtR3d05FzIF86lVzlMaskUczdVLbXsRyl4ltL7C1k3e
jLQCQQVPX1t2xiYG8rB85/LtZwl0aPatAuXE7p2eHfLRvGai3ugTqAeQVzfTa2aAEkJp9vrsvuIN
FBDTotHvGGxsgOB+wRkaqYz4gMuXBA6RgxMI6C+we7BIQNZwn4ePVJBqKxMDW+NSUpC37g9KPaVa
2jHe0c+5vm8litDjyAG71eRQVCBPlEuGQRHcbSLcms9AQBYOr+DvKg8O7A8PyFqBW8Vs9eRyYMbp
oogtQ7E/xS9GJb7Fqc41c4eQ757YBurFikvFXhoLhN8fKWjWVenHIgt8SSZ3g1nUcGOZ3kFv2tU1
usfgWX6uIyuPIZU7PcNobL0r0uCW8kwfzlI3d3mKQPbvj02LTOMpz4gGxURfITZF6e0BJJQsEK9j
Tb3jmE+aN+pV8k6dS0UcOIitTFal5TL6Yf5ZfqhmcFbBuCiiSfWwxE8gQ/gl1gqjeTgy0wgwXnhK
PvQf4NiMNZPAaCfE3CjxGk2TBtZ7GMzrtqcSPkRzU6LYlj1JOQTMiyh5DSgtVKAp+cuNRaR15Vao
twTKokHNY29hiFWPNY0syh4HhNdkXenKC0edx7lU7QflE2cBik99fngUURHVsdTXZmRvHfY4lS7I
B2zzIehnpFuJm8q6DHPorzZa9FUNq+ZWVGmnw+9dHK4mmjywavQHO+brYjgerdsnBKf2DEplq6P7
hYTU/WCJbcckyTloaRBpj7fsp3OZmeMJlSWtD+rUal4wPyeF0xUq8K/5ipJFdEwBviRT624M+i3v
c3G2id5RVc+E0kBbDZGZfy5+W6K8vDcFTULEUQfTM78TAMl95vlfyQ7Df1OksqKjhlZGRbuKV979
HegGI8cxWA5mNTQ6txPrC4N1KFN6DlfNWXe1EH1q++BU0DtoJGFRnUtA/rDQ09vF40HismTqK++m
B4zCrLW1atra1fogVjQpR0Imga12rcnObKyAOPJIc/Cv7sE2uqF7MopTDC7dNYlPt3z4GISt56wD
2YE7LbvnXhWnU7K8JVB1tapkIoajgLCj+nqTwl33tw0GOCR4tln1lIAahyLpuhqNpZ9gt9IeNrlB
HcXEn/r1OF1XIkHHkVkwMRAlT40H51DJ6YKAMlTa9HEKefyhmJg9f4VoeX+ascYBZxaC4WUfkPc4
P8OlJtTXkMmNh30fi+i/vgtCtK6RA0PcahaX0UgvH98Ll6+WOM47t0xmcFUm7amAm/+ZjuETq+JF
qDJmF35+Wzv4X0fnkQAae5EH1lNhwdD/hXpX+7cqp1ANe0Ezeyj9fQ8+FvaSl5xUuSkVBnsDMolO
zpmZG1jGYSWKcRvqLuNCVwLooxmyL9uO0dm78/3xXMHC7WZM/efncTUkoix06l3jE5cdGBIBQJug
fshobSArDvJVkeWAPWOleH9hFrlo6GjIzNd9EJL2OLv/1Y8tvubpmiaR+QgEsiQjP0cr3Q7zqW5a
a5xx+qJUwz0Iv5DI22ZT0qJ7v9YhoYxOgP6oPRgPWGQYwc3fD+FIvx0ao0pRuSPdUk8/9q3UFNYw
+HSedOcBPO6kkan6x5WcOna61AX11qIlVbucs9GK3Qg+Orys9gpHUNyX330oCxRV12OZD5J7c525
B+U5nqT55EX171YH+TV4/TSLoR9bPslR98KF9N5Rn/zPPEpgVmKx/WU5f8bNYM/ZMocd29w7Q5N8
muJljl24shM0XlfmxiOMGevhuOawuyh3FK00xe/uCWz/5xIHBJErIgOzMJn5sZ42+Q0E98GzeqWd
KQ3IXLnOH9WM1K8pulkRltiHYNnpxbXLuTxqL3PXJnvljiPEx+zeqY/u2673AbimYQMzzEC1hvXm
annuFCMgGZm+og++YNkaCDjGa2lpipM/ZUiwDB+5/eo7IGp+AuiC5VyPfg4p3FhUGDhc4I8h5oJ+
amkFsMro/kbBFWoc9AzHIaNz0k7Hn6YZ54wbTBWiektnjETtGLNLDIXZ26VwRP16gxkajzga1b1C
MLHR39FMG5J935dknDG4vMk4ysqPeLfe9cx1Ibq3VuEeUaFuhmS8O9s6bse5gqg2LtFFUuiEQb2B
Lje8ShV22XXiERJbRaZJolSmnbRC68SUOnL6KLqrA7PuxPwQlA2ms1i/PcSeiWIpg9Y3flx8ktqO
SkBOluabzzyTdwprsYuuueaRoc73egv6G+jmLRF5i2BjiQE19kq7i8n0GDGOedmg+iHHKDEQJkAu
GjAOT2IKH1U8DpVj7Ynx61E1OjKrPC403hb7lL6ZZfNYJCmEnG/bLZCR/pV4vfezvZaAIjp/vcPp
YgsVtTrGzREp+QpgMScB2YdC0IcVahnJDkwtRD9x4omeBQ+bs4xMvrKWRVNNIp8QflsM0NcfzHHw
XEF6Wx4vvDjqq0WVoAUGjZ/6i5MdPg19ptLOP84zM8rfmhEVLnoyQcWjGPkZoyGhV/SYXH70MiDB
78ps/xtBGQyDEa9/1TDgqXNb10toL9yfXX122mGcMqbXdaJqsu16kf8hYQF3o58t+lmXxHMoq8r7
vnAB3V1xU3JQHzv1gh1PmaQZnyeD0ORFS0Kcxz/5XmSt38f2SIPcEkeJGRklekhvonBJluW9kS9W
ew+nGYrNjpQuu7TXYYrIZQ1ApRBGxwkhElOL1iA51gqZpUb4dwAbweg9rZ9kKoP+rS6rD5eDk5dL
M33NFXMQoRdITEM8nspIeTFeANvzU1KSVf72NsYZX2+Nva8MflvRM9kwBBYmh5LeN7wePEtJ3W7M
/1i/l0hwkIxUi7CILp2LTk4NQyrIVmX8yM/sy9w1VplSKa+wPBexVoQ9oYdKrxSuPu8fQfcDoIGK
slsPVOsf/W4yczJg/zUNtZHt8Fp2WP5CNZrmW6vbuiUbtmAKZRv1wl+/dCnqtZoTWjH2KvjUv4MJ
k0ogSW7+XYcVVk6ylD/9EgWEqVDn92uQyZaqepFJbM4fQ9+MKNq33ycyqYdsEkKM2+MqyVrj8v9h
KPuRiSdSovP6tAHQBYX8Dnd6Fw+a60WbM9N+C/7pNxydlUNQXOYCELpaFwxSACqZLBdGvxO1EToP
s82PpNnLChQ2hFJuIwACG6wu84XcUtXuMH5t400lpEieNH6b/vMZYm0kFuEwzwPz/GuUQkDZo02t
ZeuhLeqPUfNfOyK+h9iz5UHNNBbWuCExz9YkpoE2fOk2H+lNMW8S1MJ4gM+sHV0m4+r0jrz6sIld
RYFOkzUYSakr7oOL4dc7D4DKgo/YvOCNz3exFwCAOWmAPFq0AEOM+xWIFSv6neCFpMnmdy3Mvvrz
TRDkSTr/ANKM1neWKvVL3hEHZ8P2eoAyn9pZ1tl+p2LWee+SUiVB0+BmVpq47M14q7MZOa589PaO
WQ0TFzw25S7GBuL5VHqkmxzO43aaZ5EUC8EQJYdvO+JfuTBvtIVjG91Y19JYk730eHkn3A+SbHJ5
zJBJsO5y/9VvD410vdC1908V2zx17+6Z7UUnLRPUfkWM8lvJOXUsSzwxP53YDqwNha2MmIG4E1b4
/zENizt3lS+f8rhavM4NrbQzrP2QQBS1NdbX+RUmNJwujuJ9+Y5OH+GdmVEekM+Mu+67TJ/wD7A0
qAc9wrQmkLVQYvKRipoE53kTRYGVzxlwe+L7FLBfw1baiPzdfXEF2iERnXFM/SzeDLZE4YHEsRf8
rCy6Hq/Uby2sIF27fbY33DNNmPWXMgsNMdYMPGCpPcf2cMqzpffwvTj60DDJ+8ebJ/4i+RglFZIt
HFbVtYqSQiBMvOBYWpfpoIDXm5q0yRe9iVl8s644Yu0cr2ZjWT7r3M6xdtmHT9Y9DYonymEry4Z9
AA9FAU3TLhfaxRlIQwfQaj7LvcIhIsXZwdVjTknW4eulHM2cQlgs43TG5Hp5eKNFne8TEJn6l3Vh
qFDguTtYP8g4SmdKG7nhyQsLutyypRLk2G+NhlT5P4kSuYJ0GWa+XF4lgjokM/LD3F2SgpK6aLEC
EjrpVSWmwvRp9LKzl9x5HVMJhVX5We7zpLTEzg4Q8+snZsDKEk3W+2DKrrn2dYAhg1qnXqyXOpwy
vG4QWjEMapaUu6jd7RelvsIe/CVs/RQpm7cWv0pOJWd+170V24Qmj2sOJ4T2+mRJc4tcTzIhMRBw
87VLXc9Qa/ao4L5foZaxemaz4SPSZpLWogk5INKxgjCaTWI+k00VlqL/9X7MXiuyz36KVKMYToV5
5f2aC4lb8JRk1rxB8hBYSdK7UdUjfhcvbcEDhnmK3xrPUOsEf9+LzSTU15eG98eG/uK55z8LCMtI
fp0lEA93gJ7J8C8aYfNHIfAhgZ4k/s0bMEKSCpg5RZWVNJrRMYJeJRL42VVCO0LCFncjdhp5Olm1
M3dPPmuw2C6GYskYj/qWhlp55I0pSKDK3zdU6Vwd+bV4F0hzfUVYsJtyuU4wKjxCdIi4APVyCTZ5
Y+s/GbqTB+dDWwWjiHTSa6MIFBN6zHy8MZ3WYx3icUobf1DTWZr3T3LYpfoc147ZVyhfMbQgEufG
7P0umyLf5Inj83pfQ8/ADWQBQqqh4LTLX4mSR4qkuJKn3B0NCfD1y4SIQkeL34LxChwCa5UVtOB7
9e+6HPCZqbedzF0OxpK/dIyisZ/wMu322Nx4ytu/qhFJ6p4TNkOX+OMedsfSMtvLzKTZRn/k74m+
a0sAyBlWqyVLIVbsAt85Xdvo08zBed/wl0vUqdbdwHi4xQnE43lxpKALaztLHUN8xKHvqs4LuT9E
sa9e5Ko01+IuMg09QOFOYT1E/cFkHf68ywbkV35hG9EGJR2tpJupKp3cngVQbpQC3tfPveBdXLEt
n7KWC7UzAJuhARVbB57ozn/XkOv826j49TfZMFF4m5yFw85D90S206duVpy+BpCGTfBlcw9fzyEr
Tdzwdwz/GBBoI5GxmM7tTrSxbBb3YG3t4sHrJa1DpC/+nHEmI9cRbXNroou1rJSsCxqeXkvcXtw4
j/u1qtcmfqxQo0SkLq11Mh7ENRVPcS0VNn2fwHgQqyWrTRr4+HOism8VYmdJza8L7uu19Wxtem+P
pNbu7vkGJtZniCuyAgc6yhpZpd0XnKEd4GFlauFvbMHJyY2RJjcm6TEj2CzVEBmmpbx50CTzZ5fP
tzY4wV9LcD9yCMI4ZLt4ZUvjC8PruuiLqdNLKtjOwtQ/YtwjLJUBA6cUlVr7I2LsNzJ8tz5C8iaX
rl5njTDIapNlKNY7PD93Z0CpNyswD1NvAcomiQp1AVwGPX6zPptmiEUBvjB3VeU+EeOwAbFCnNTu
6+B9nxtr0op9ILOBBBoydHXa2I1yScfOMr5ikRXfTdK2bkiPTjGPyq7edFJkJYDp8tI0nngUbpnv
Md4lw6KR66BbSsTduk9lfSIb69HbIto0Vz/LsGjHcIuZsNUYEonv2TY3pR37mCl7kDaKSeOE4ERW
aAx9XKyI5RbVYaQMGTGq605Y3aL/1yJQ4UNbqgi+An5G007zvhCPuG7WX5V9u3CTNuGF9iqII6Ll
IdKqZedPoeBJJimTHfDcl09uwllV2DQKZ03RzxPyjr2P9J78iawcKupNm3bzbIGUz1OqThpAELgK
WqyYo4fuDquEk600/peZ6hwgBo3GTcRQTwTLTifOxtPnDwg3QDUTux6NOzG0i4RkmyRFN0cDkBM+
joXeR9zeE5InYVe/83r6kaTzNclVPRvkmNFCjkllMl4GC8HMYu00IjJHNonuNvjibRaS/P2ybdaL
zAoPhStsgylt5JLVjH/elnc8KVyHkiJ273P5MR0ptuEucscvMShNcwitpgoKXEKNLynLsE4VrVHH
HpDO/unMi2xI3x+hsqCkmNE9iYW/qpwkMuXLRRhPv/uXgUXdE0psEAS6IWUnkQ4hD2N/aq3nLSlm
OqKIkAUlbkd84jPkdZKiI0OjjEFU9lzSSXDjhu+py+lelyDTq6KPeUDxCBpEMotpcGiapxE9UQ1u
j2dez9bcTGNZJYbZIt4TC02OZNOsvwSItdMKrmmYdOZGWLaZZG02CrIQBdcFaNLmaYiMQQdOSE2w
s5cu7aOgmeFk/D4AqqDp1gYn6CaOXc5qFPi2s8cMcROXnTJdSXhlVeG0Kth2iv7YLz7dSucC+XST
nJDJqTqGf3csN6ySBr2Cf40iCClmbmvyvDLw0eEZnFKWvXYn4zy8kO4gw9sK07L3bsprs35J8WEX
pq1hcRn6oeRdkOYqk17HhLZ7WxZdBenm19qjimKL3tZQlTMaxxYJ+P0LL1BdBu0fFGD1PHZaI1uQ
SL9JMog9KZHDKzYghw/sgdc5g6FdvoPGFp7whiXGx+ILyNO4CZpyylza1JahJQQQtZ0abLHOiLZl
feByJvCgRid37cdJ5UIFF7+5NtJ0YUN3hLCwmGyqC/AQowT7pB9K0C8+FAS5iHgCxCR/KLGg4/hz
D5rxBvGWxP+S8iH13SngzaqIBXnGmpW6UVXzU3smQ9WDAfO+tbQakmoMKGTEXtehot3FiGTHb285
363uecgJRFR6AVG7SPbV6mnOu50r0RT4h9bqQs0gfw65fyfXX9VRugX7SFtN9iBS1dYw/riA/40X
MQFs1Ef9ldB2G4MgO7Llfaf7Ic0ernboo8Bg1yLWDciyudNFzL4zUFrQB0drIkZlg43PazBvXmLq
sMKyZqp30LJDGFs/mIB0ZyxSqQA1ifkWqicMF2RVyHvrUYayyyJEl10944YxdpfWuhIZ7TSaQrS9
eo/9TdYUBisr99RJMWUoURjzc/QHcB2mVMg0TZPgwi9wF6cgwQenj9K0Z192fUtortE3U4FBv705
y7dzhgaQmodv42FBBuaJ5w7YYFP1MffDVNYePwkBdWB/rhDZZljDkk7SN6tvZfnVwgs1u0uQ/Jx+
z4g7gWm55z5COwbSNUQVgKufOi/UddN+4abIjJ5eCYmcAxQly9M/nZSryeucjSZL9KgJyqUxD60x
yd4Tjq5zLOt6qBkk+AYwnyHnTF3yYR7BM8HBzAhQfkFu0UfgKR4i1f/9tgQMNxnPq0oTcjHmRwLp
IHJqxn7L2W7dbmtzPHoWVHwcfFKGeAteTJQlfO4ldkdb571BpEdQGLFzWFlAv2kNZ45fxM6v0w4R
VI68E2EJXqtT839GDVauS0DDerw7d1k5MH//cDHn/0z8Ql0TCPdE2No1WIjIzr/GxP9df24RNUON
btqIp2pQRrGMQphwD3niC4PNqmCbeU2lLDSaoqLH3iu3nDburtQjjM77FjBuE+StcNRCKFxmj7BJ
WyyHLS2vFIdLn7KTQfjhDtKdQUauVKypg3TNMGryHui2CzDszJFsyp8XvXT3KfruE5HtrKtjRp4l
ZuzFOlKHY45PtkDoDTXLipSLiDjchuZQoTbdagLV8sAkhobomtQu9tk/e4Bkj+EGqE421GyTVerh
FJLon/4E/JZ2v0SbGOw3Tc5uWGOtvqKpaKNz0sDypTahWbmpCdm3x0IPgat0Yfa1zq/MOx9teTHF
ShCW8V0LX5gz9pyrXHC89nvVhzoilPS7iPOi8Clef+2q6WVS2Xtud4JA5h+sqxpkNflP6EoBxl/P
G2+Pq2yo5zctxvPqNIJkO60VRMpxlzvsSrfxTA1fCPCtIaBaBY4E4GrjGvosUzZd8kQsD1uYEHYg
HHcPYXMezOKTeSoheQSpwKttfdolDlv4ZXgc7KZzhm/56XMjfFE2omwaSz36Lg2kj+wkurWmvTJN
2BGwUTuLdkOENVC+uW+mN9M8l2xw2hZ1aHo9U/ixyIZGKNtrTOut3sBtMJLnSfQ+6p5j6qfuSjP3
iV9rimsQN3PbiQXsZgU32VRrNHZdUVHUATFkxcQX24nO9SkXMABUuQa4vS2ZkADJomXQNcDKgUXN
dpA0iAXJQbwkPGhC6X8rCSCcVW2PZZDJWqPO5RZx71e5QwtrOQTBv85Yleuqjq2xbf6+JNoC1zLC
iZbYviOlAX2Q3qNOCl/9SA+4eA2Jmp7mJ2pafY2S7NmGfbzbaxQlYKT3JShtNknNwUSKuyv/ELzQ
oYXBeHYIAE8U3UDgAaQTNzKiAoAXKni5WsM0mUGeIJh/9BHZRKBF93Kq2vqsmKgEGpG9hi024UK9
lnjWcVGfqgL+xa7lGkraGQpJZRkcEjuiiZiQI8rq4K+haxFz5N0Vp9YmR+VKevun8EsaPNPdNChG
yb0jACfXIqBKKA/chdGqv3EhGsN6PggVDruRCj658swXd9RckatuY4OLCIWbBL00tlwqETkLABTZ
CLa8dU29zQImZlyUEIP3XVsUCo9l2l4QYvaJmGYHZAmDnfdz5RCB10fziX27118xYJdQcXTlGsbE
nondiWdaAoLg/EQtwFCMEVof8sokrSdXts7v4K4hSjkgjAHUtqHTylG8eaMtLkJnpyNPtuIIIdYm
VhhU4yDsXp2bj5BquXLkCVD46ULcYBtlEZIBa7NIM8aks7EtFnUfXEe6B0qxJUnSdvcqhxRKfY9r
Tc2R7EKo2sr8uFgH+uJuJ4xe9cRW941MccnuKLn28XC0po6hXHla0Nq4ELYTri3U71A/VKII2kvb
zJCyPoL+1BllB8d1Ir2h+CfM/YdNKv8BMWZd+JLs5UKjGwkscR15+Ad/TuB7ach6vvjAn0l5GI/k
SbuaJq3JAB12owIJlSjQIzXptGwZ5EZ3FrhfBX3M0TJuktKQwNTftjTzUWS+wZWP1f9uBgs9LDMO
ZujKiJFuHnghbPXrYIuNlToN37FHlamKn5E2CsLOgy8KhNQkb2XGKa+nOd+7ICREYyKwpzSHJIW6
jaIWN3eTg0etqEbF2Lr6yPxSLDSsKEsW1/8/UGAv3lsp+g9D1theUfXV003uS3RMSW+llLtKzI8s
U0lfr31pbTC8bQK+MGUFJShABBx8VvR2SRWnFSStkNiK+AS78fze06PNT6G/rZo1w6kwVnBnwtxm
mXtwKQxmNL/IGefX60DjMXqH5e5Dz5R5wjU3QWoBD3WAU7WOd/IyOtA0VDYoYiKjwUOuoW1sG0BK
hgQtkw3WEIBdylUk0/MwewoKXAwh8NQpyqvF4D3ObcdlxbNlkna/1mEmG700UvJ3W69yGNlxI+h2
y+Y08cLT/ACnDTXlX2Z9hh61FC15DeYSTxEcLYnlP+jWbm2de8YfNYwFq7I0BqGPf4iFiSIUFCvY
sH8KzbdCD3lUfPDDNlQ3Dk3ujio3mNJX93xrrsxmE9ujPkozHXKf9tz24Avvdl5Up0EIodDc5L5F
O6Uwf6M/+TFYkce2XCxeNFTN4bG/Ez3bOLLcAl3Kv2MltExXMzr4QO+Ccqp/ZglTtAcxiiC7/i4m
oEmP276EHxdFgR+FdYApX+tdiCuB4GwZ9QdyCL756HWroSdSDnVktusAEVhYR/F1XyTK7hBmvmdb
JbAmksVFdz3txCbxg8Z4U2KETEVuzqLlcXgYgDqiVFLbiPaIX+TvRpD58dwnp+DWkWH1Ec8QoUZR
9LGNJT1S8+lb2eh1cXUqXTcKvsiySp3n49MSuffWzPU8K9GsqV9cEKSvvE1nO/Z5z9cttJpbQBZv
oGbmX3qKlGmSXfo1GR/x2OjUIHXHOQ77ECCom4HrTRykA3E4ph6XvCOc0d0I4Y3Uczr1EDJT2Sge
ZA+1dfwEObQcmNmIeO74qJLlreaZ0cQRwCQmeHYW/8DERv6Ko8f+Q63VdcWWFe3alx1WR/AkHSxn
xbY2bmT1z35m9W1UZTo7Ed9gRY3xUsUoxoLw2SO+lVvUj0l/UXI02VyfZYz9Hb/VUbCHt7U1ohY/
mbLxVKGf9jTzWBMMzT/TQHsQyK0EM+IbToPpz3gKLEisCZVFDPeC6lzAZUWQV0bSTCcmt3IDPYrb
a1hGbIJEnuPGitnU0eZ/yvXdfnzwikqiSZZFAXGuM0hQZw2ksWcIS4Z7114Oq7DdcRmd+4qk2pPn
PWkJd/lSb89mlHL+EBNRLWC809qCpDNplHEOuUkS8X6eYDMsapx7C/lx9Rrs6fgyoaTKG+VsIavF
JiRC4wAmoA0Lqh5vVSdBhizu541nLLoXIUIcCmbE1IceoOHLjhk0foHOUStepN/Z2w7U6hYcJ6Vg
3gyBxRBX5E9XhwwmFp2OWdHld/zFxcY2u1U6ZKIZ0XpFlC2aX/SHZLf+KS/YJlLPsU99cWaW24sx
KjjcjlksTZHbwixxaw34unT9DoSnhtR7leR4RtqVYami/6JBBcOyakduX6QS3eHAthZCdYWkMKvw
B439nKztuw5jQ1/heNrwBEmLJf6MLHdNe5mbTxiUg1kqTkNtSh03VhTbdPlLJ1M3sb9WC/7ABYj4
Nbx3Fs+SbSskXHZxz/oeiusUxnKEaEs8FLU2tUw1GQzDETQ7brIOzbJzbOgK2qDrN5kz5v/hGSrF
uzl3iLPT5yN8+lcYiqQq2RgBjKF4E/Q2MairrSO97lXmdI/6UFbTtBnznOHnoRwUzD+2VHVGZOYB
Ar/j9Eq/sBna9+x/POjRKRlZNXvJtcqsz5XO7FgMBy7jLEkNkMTTsoOxHtskjmoQ9Ymabzvfp7Pp
GxCA4OVa6FcAFI5Hy264krlVWsIj1APPuz4l+xC4EkzjUdvE8d6/hDyoVAxxr+1A2A4GD0YxUEd5
um66Usm2DwbUX+or8wTluGCJXhRYE7Y4SYw2tPz/I3UF2i9p27lx2WwkePz8zjv+4WtMidQ1GRq+
dpiFX3xjLwF+aYXzMHph4sWy82kYCNzjFHskr4xQjzSYOE4kWctsREM1j9Dq93lPcmsvzGgpte9H
wQOlBz/v5wzcBgwzMI8ZCtzR4668NDQSMl1OMwegayv0DxK6wPby5sev4r3fKFUULFGw4PMmbyO2
5kmiObXWIrxBbLMyToxr2WjMVi230J8wz4EMjVAgtNd+AFGQdVcpbUjqfx8cQSqk/Seq9jp19bgn
hMc5nVx+Cf7duP9W9Znmd4VwT01b0AgokGrUzVGuUoUYTGUI32bqkCkvUkfxEZgyKUeUmh0UL0WP
VWkA9xfiXDacJUFkSJCGZc8NVwoX/Y1hxcMiQKi065L6On/YLrL2Zj3RA4wegNNOFl8NT0blmek3
k7fdvYSd2Vj7HtUCel1CGnJ3Lw7Ub20jVzX0porFadFPRy56W0oRCtZ9Ry0vD5Phi3zqSVH0MIb9
No+eawxARPZTUCYS2mom6FRSLjskZyqXOw10TAs9c5TsufCKrCs9ZrpNXskMdqRSBu5vs6R4WfHd
O5+6pxzfg7DgqciyZrcgFjWTDcocfnita+1IdpiRfRqm03ATxloU4cF+r+L7sGg0Xb6CrJf0Py80
nbdWZ2Wj1U+x2dS1LPB+Jb5VZMYcpoNTr2kscdY8It++rojBkPvA4gmpmSAxTXnkpyC6b+VpOcg7
yfyc1A4p2/AJD+Xb1qglbQYTp85bNSlImnZh0onx8mO4ofJP2+B8cUhihtn4Xv6tsvipkAUXN0ed
zwVSczAIvAqpMUgkodt2HfpCjZkRxNOp41CoaYJ2XIYXfS2+jDg+GlNtiIk9sRgoUR5HR+KSsmAU
G3Vf5VRJVqjFRXRzE3KjvOXUSZaHg1y/aj5lxS6O1XWJgKGA8yLnnAVjgL+zr5R7va6jpnLOX7kC
4IaJ7+8lU3vx/XUOBMP5IDl1AeuY0jle34uP6P3xw/MQa0qKQJElUTP9bNsKR/rbcuugvw4g5UuA
uBrl/sNTHe5lEYmq06Sb+XogONWfLuhF26LJ1Ap129ia/MGX7cawHP9gDqf8hwdziUCrJ6r2BVXk
Z0mejQLaNHbK8+2NzGL3jqeHXQSSQfDvlDnQPPVslS8StzHciGRZHz73Y8hR4WxgGHKahN89DBlr
n43tKLy6okGXE/G7dIVm1clyu74xUOQTGp8dZn7b6s9ziikW+ho6JvQDxlMCWMjUuX+QwSpe203n
trewjymaFRpciCuVfCRM8ejgBGx5wBr1GniddC/2S1H0OZ94NgBOiR2gAhFt3ZpffQjscyAmRxRM
Y3KkMBwzhdpc0qaWrazUKp1Vy4HKu348a2XZDpOBlaFTmbrYNc3m0Pit7IB0IDmLf1j8a7mLUfbp
yeXPGJso6paEmT4JlmJOaEsQrmeS7ViJEJ290VWZbPY6qLPP+D7x/soyiyvUdbSWCPyFITiMkeIy
KcDvqLG+w++dEr59FT6OuHhlai+R6XI6SgLKjO25Sd2//cf5xR3sE+0P4/C3puWpQ+uC5yfLGZdE
Xs76W/qjKLo8H6zd3FZ/fF6QsL/jELT5x7szH9r47dTWfypW2nbNPflGPYhPPWOuyupM6DB40vwo
PKf3OntSgh8VWn6rJcSYA/2Z6kG7CXJCr6UYrL4cCG4sPefjgi9T1nY5606qNHFuCIrAfrMoEPU2
XsKzKJynAtrTlPS5nwa3a7XAGq34HPJYs1Xqj/siYaFFKd1ReXAiEeKoHjTmLp6A5AxBUuv0Us1O
wH8EOdVeOSXeEhmzNy/+J5UoVLPL/G20T/pQ/j0h3PgMCt+naO4mRB0RnY4dQg8U0kvSL6ETiMB7
hJIvCX3Ai+xpWy18aixbAyq2/VTMUnO3kQtHgWXY9VGmxj81uOe2rgCht6OvOHUDQIjeVTWNL9HB
qUeIer8EiftHY/FMN/Jwy4G1h57CXA7UGlMVL80CzCkAxQilYppSZdVg70FV+GEIqf+Meyc5e7zX
11HIps+MIuJKFSdXmM+38l/qLZwwJOVOX756K/ndH3blkV656LJXBOVtO6eKdDEfQDo+wNO8KHwb
GHj/l6zN7oF0R++zVnef4Mcu2nb5jbgC9eRsrCH95TrT7VY37soZedFkIapCEoEaNTs0zfuT7/gu
4YLVpmh5+IRIJaNhlMPwiMERWhovJxu9eFy8bvXz6jyuVqPehj+Q4ch08PHYul3SAACUffZsQTz/
ZxsQ0Rgo/JH0jUOx6X3842u2sIkNLOpYPjmSavpmVI8f1shkkzKEogDcqMkreq94f2atuoLRC3OB
XVatcxCzwEcUhaV6mlDNmxQd9ksZWr756RjOOFQ4z7SAzQnpZ0dU9ZVCw0iaTIaowOPmi6LFriim
jVCqbVKNORtpv/eEBhpsy61ISCJEkRx3MHtBBtkF0TzwhZdsk/L5VW0h7lmLi/a/MYuN6OCYdMV1
xN5J0sJJo3JGZ8YiTg0LN2jr66g9+rLpsxAO2QO15ExSYRBO6P68h4+KhCrIgNGLZ0Ezkp54FTOc
6ThrNRGdNtOPoF5sa4Xk6rSMVYAYd8XSdiGZPUYHF+SdWqpie9vyjCzMJ7WcDK7Utt21qj3weyzg
J5FwiTRy+otRW7G6YNSG1UjWdo2hS7LD32LzUd89Vie2zRyaP7Z8oe7MuuhVeYWMM8fg7bfkS+u8
JrLLxvux5El4aOUHvRypmgBBUGtZ1+WjqcwESEunW1hNInF4akByIod44Y9rq4lxAmElTnD0Duy+
vZArbSxaZIRFUVHZTEycXE0/PGZ0jUm1YIFN0pp8MGwb/n2fZrMKLbYquLP9zgxxhJcHpaAokW/M
jEHo7ZUogRF+hXjkdvFQkDgbtQFrpsZcb8ogYLHC5dIP3tT75JOk8r/8qaFmU/le8Uxk4/G8bU3K
EPIRrg/1oVy9FKONoCqWFnCQik+s8BBCETXBplwCp1UAF9J9YFIgUgciAqMwRrTEu/LJBE4Eb+il
XanVgba1QfGJrVREijga4kjp4KnDVBRL1zCzvqfEsZFlR8z7Ix7ghg4NpJZuoDX0lUrBjNMM1BgB
O8g6qborW9u57DbTaMvIJEVtBXCGpU2Wh0JXOqJwdHrSrRjkLF8ifZ2ZH5ATWDOkD5L37GwTwTU9
qQ6jaVA78KgunVIqzZPqsKp2l89r+1ZVwkHWMogf7Pqlb2irvSa5dL/zmC6Im74DsDgfx5BUTWQB
lIp4y4cu/y7dELMEpWuBPlWXD92UWzPjdYpl8Z//unZhj9AcLNQh/L+gT2TmmsW1k6XGNwJjnJsk
LpFvDdfwznQm6HUKZ64MnToxdfVBVjrNQVxOilOCXw9heVWCrzpP/K8JJ3Y0BR85fKKMoRUiWWbn
sVCLkj6dvG20SssQroCyg9C8cmFArzKkkNxxGevbYwywovESzkZGfdi9e9UmFtYd3aS3T7tUbktc
6EQlU1m1qGAGolN7d6P29fVCviduRmob2fr3AZ53dBg1FCJPmzRr5ilVkJtg+v9OgIteVuVyEvpn
fxkyEi/ECNdke5m513xcHAgdN4uMdh52x/kKH2xDyEtHkD76sOx+KZaXo4LJoH/AA/YW7OJkeYGN
jckXKF9XviAMtf3iUG07nM0zYgJ8wAeMcekb7t11rdSa8W1IF/EI20OjarsWIbx4EyYhbiLMTu2u
RpffduWY8KA53e87B3YOeERrr33JGuZqpYrJJH2nHzJw2ag8EIqjr38USCQrz0cPubfJogEXSoew
Ku5cFPzKrIbGT4W4QUQ8768RHIqr9sBylLaDeJ/zriSigBenAqpVU29Mo8TD9v2TlgV5MFIeI3hw
gHVKkJtG+uj3iHXnnCZajm0OODLbn+BO0sj/irF48DlM2nEg/gP3UBI2pt/2YqTvucZaRGqAdtFG
F139BUaaC8zMVz6buCyzRVGFHlTJSMqa5F1TPO/zD5MoO6CHPF+XMAxPY84PL1jVh1YhCOuv8//K
PnixEee5xd+pvPKOwdrfDl9NOBY0N+7qTsMNGnJp53wCygfq8XDNLyZRwV4Jf8YAiSej+M/W7yi+
ej/uKF2LaUvGrCkSl6C4punlq67CZBih0GcaSVrdBYMh82Z/pAa+nTC5ik3W2krwdZkmyl/Y1pNV
7nLgQ5V3ELjqA6WE8fKRF4y1YYeybOePzBwo7zUg9sQSkYKVAQ+W3Cqb1hGQ23ea914Ks5knpm7l
OgDaNxZx1Pq7neualy+tTew9alYH+U54iG3yMg5UkqgzrQwoaBJJK4SgkozMYinGe+86AKUmnlAK
4rO7PYg13U09fkk/8zcuChbScoR69/NuaCoa3K2uJqEkQFLODPGZcpmQoim8Pd5SEBRh5Y1LBDyx
1r8nQ5d/vcBEam0QkbSTUJ7JyCtoS0Y0Xag7lhmYqgslbVjuYds8H7H+LBdxihspZ9ZkpIYNN+l0
UNr8rmOjS1MxddG4L20NmB4uRI0YlU4T6bUIAH95jromPSgCuAiQI7U7AmPyT7FK24dWJ0wMpSAr
Z9o2qzEV/t1VhjpwvOykS+KAstteQ9Sp3PIQ7PHKLNNr/QuUWwJhMpd58EGWK9BizL2z5Xnzx1gc
5VFw1Nz4fZzHwo78xngxrzd/XJ+zc+dVuZ/BJlc8rHkrIz6VgYenvQHC4BRn6wp6R3ev2fOkCdCV
VRtSUICa0aGY89SxNVuPlIZr8c1Vt0Js1+UoJ4WshkE2SqwCRS6vwBPwZHjupOTGo878zk6RI9oI
/YMXvNkWOc16RYoPE/WBGZQUwDxhi0IG+jRIa5s07fjIYlHk9O/WWTT+iavch310sE+XjBcobIZi
Eg0s8ee/iMxssc14gWIorejEi0jvzcT70D/p7y2ApugqNgcEpZQ2o53oDJ74bFG5o7n8JY3KCJUK
5cxfPwM0fdDWnDn864W92I0306UwR1YccqShtBcModgnZymWyvCIaz1rl+JsJ97o30EH9TGWEbnX
dnCE0S/lvCRKIfNidyoHXA/6qu9zI1GYj4kKR99fGC37aAs6uhEU94FHvtIEQCSJ2g+2ZsUXw8aP
P6c7KwgpH4e7LhK0Uu8Na98GZFjaF0QS7KO1abMv48iOnLUNLOvFoPupeASPlmbyJk0b3GmtK/YL
+4+w7LDGFfj9rOwTq1F1auh5jyP8UnFkTb8RNeKeojkUckyfCu02SkksR/KxH6rcdLlNuLCOWfco
0+1dta5I1c1H1qDSWQ+O7kzNL+zltVdx0Euq0SyMssMf9DK0ixydY5tdRsxgufRTDNVvpA8+6RVK
ChrRaB7VyfPjujRvHx37euKTQ+8hMQddZr3cplIWPgAmD7EQ9Aij6cfIrs9K9A1BbaNdKZBoDtgK
L1EzBroEhqA742u/Hi4thovSeQIZQJ2WiYawq6g79MVFnPfwMf9gSZRUH8nIrvoaIli2LVIbJ4vW
FLSwX/WbdBGC778NmQP2E5/ft4c2166bH5sqrO+mMFO6U/KfsEAauIahniDfEw4h9xE66DFOdpm2
C93f6OfcRioufMR9yqVDlH3r8rxXv1f8idtIhVAbi93EqoPEiel/uua1ielez2DHGKM0aJyNYZdY
L3tv3rpSP2574HEXiAmDcLGVjRaTSGHm1UFjYkxDZNxb1M1lmHsJKwMzuv/awlCpJ/Z7+MZrK9fs
aIDfy9hoM6vwNAWl46D0PwJxbyADTDVpA2PSOyJun6L7chvGHVuAiFnVFozMg0epPIQ3wHJiK8yd
Q51MXXBd3KOnHs8/9C69qiBphK+FMd/Uba0PNNvIcOSB2cdrTumvyLYt3lw6UipbgjD8iHrFAdm6
nwOJ3iRElPgpogTrHjGgsVuDXX2k2Bw8Sr7u8wNBthFNXLuiJl9X8DWruWKasUbPa2dwlfuK/MYb
sKIK6UZrrrDIeUdgJVyi97xF9w6hWnaQ5PuV+ChTZWsm2MpaOGWumJ2Y3vbRM2MbrhyAY/p0pgs2
1NGiI60NzuF29aba92pqFGVh+0m5JycfIdADw3X31+T+/AbCA/WWIJ9tTUqb0ga57ji6YoQr9Ia7
WVMFoEfB7f3xHNJL63UBLAu7T/K5IsOO14BGQE4yTpeCr8YsfHV12pD69prrCJQmAro37erPlwYX
x3SGuER33Mf4gwA2wusX26ykva9TljXb0X5+S8pWxhyuPoV2H3qsGNbSkiRO73Sh0PHi3NARg6di
mjVoyPiH22qjmGR3NJ5YTJvSWlG33nyK9glVTRdkH+Idb4zOLGv58kKPZaPcdXGwc29rZP1thZsM
N7qMdX3prJ5z0adbCpk8E/TB2fOZKjVA3iesGqU5thQaX2ibIi6272dym/XMCaOIxc3pVa2RVlUI
oaX7eRLrqWIY6PYVDXp3lrh47aL8iLNCSwQhfzM6f7mtAcdv5Uz33efMjkoiww0zqg5hXrqIaPKx
w9jLc2yagceDnRC/eS09wkz3P4VzKJ//hF9fqHNMtp5XHwzGOE0QF8o6BWh8hcCMW2Qq2ZLnfXY4
tI1We0bAJzK49GWxYbyCkoiAbNHS0SCrC3zd3deRDwIanbbCpBJg6BLQTwZ9TkwHo/ODQmSxz9pY
XLxVP9cKTEa3I23fIfe4jnA1v7wjjWUGYO1zKweCx3BpvR3Ckb5vPXWdHu5gEM9N0Tg3waj8QF2p
tdNAZpGmQjfm9nWgBYAEq5Z9VE6daBLuONqA2G8oOLR213NRweXFOrSTLs2W2KEGbzBWya4QxpZt
y7B7i6rINtPlawS5ghpc7/bhFuqw4NS3WKTmPzYqNjMDqlLx4fgVVp9gXQaxmZsGeScSrn08GDnC
sRXENa01VA1ZcPdV3QpCASwdfSP9Izu0FhrfaEObZH9/mVm5oHlmc27Kzo808GzACFl+tFdm/IjT
CdTKuyJwBEqNSo9gE+DhtDEkZm5qQryP6Dd6AA9SBN0/uVHJ68oX9Ctl6C+czIHWH1XOrzZK7pZl
VRSrdZbCQrgy743LigNwHguBoS6atUtk8julesu37yd97W7E+n/P24Ymwvk6h3k4shobl4dYQ12J
lFS0IZKYGpvwuTN7W0ovBLeKUZcB7bJ+hcoinzSXGJtZX74w44m6cMLjoouGRs51oK+3VJmGzm7p
ASneq/0ZNyIIIV/kMd7IF4RuUS9lZ7NbVAVHA6idGjOjKnDa8o463Jvyc4qq9warWlQRG+6Huv5l
s31YVBuYPAAr0d2uSZPleoQqbQe5drJsx5/n3ah42zDmbaMLaj51j+Wep32djLALtvnFpE5edwTG
aALs38tCgy9UbUmNmneChPWJMnjaHqyU4UM54cStVjj0+Wbqhc3t90BB417Wp4R0EH9lXuCRYCEH
OMzR8HSQ0cva0kPhwmrT+L/GnwEFvgzkbe3grdhDUJik+1o20+Jq5ri9ljyI7JFtV9tfy7H1kJO9
j2j3vW05BzFPpND26OQ1qCxdldom6znJJ+a8gizfTE621kQdfeIG+FoiGGNqkBdpI+LcQt9A1Z2G
/wSQTO8W3Es4+0FNH0wdeMUvvU9oYfFIi1ol5FRm7zZqLTNkI/Lnrhdk052Hr45bMIBcwhe9ySnR
y4SYwWNykiiBH90Lz65i+Ws6uoIAsH2FvDyBHuJGl5i0iJgnA2KdqkytVeUl5aOivexoSPag1AEj
fCdl2HTxq6ktXoZbMsO3ghp13znNanejZsNTFIpB1KxUknZpUy26qCgjmJAHBoXlCFG9NyshusuD
3zxzuiEfheEavfYTowkAJHPhxzbZouhOjR+ueILbZub0adGoSpWKyWBe6s7VtzCtW+4/KM11nzOE
kqFXWZY1ivB6qJVOSlhUo5zPzhiHBJOKQWX0YPMrI2ODf/o7+BCA4hqtZMLtu2PyETkdO6GmPPa5
QJVKP00PCa3VYlKbYpHoqaPSSXLZBPjcd5/LPzA5nsLG3ZitA4QARw17LOcW7fbV+vOo6MHu6exg
Jx+Bek0ZPzJKnT2hxmqknnwi+v0yS30VUJkK/ySj0V01vvF3vkBum/7HxjPAPXVOvm9cQcU5LMT3
46KGhqCOMM9d+KkM3AbuNKe+cYpboI869zsP87rBHADUbZbm8BW4DfKWOhx2/UNVZcxWQnIJXoI+
ht6PTqWgs1jWBWap/KBBEi4Zm8Yz0H2jz6Q4MNcjxZ5OQuzraRrC3PmiT/3jrvdIU+7wa4T+1lDv
QG/kz974BKT3/8AJ5LkNrcYU4HbGhh5GBPCI1mocOP0MYVuRU+zmi17AT3G84elNDSY2HmI6SXu2
jQWykvs/0Rw7jWyyijGXCw+v54jwiciKsWJtNgjOP/0wOJ1Rd1B77V5gevt6gsUssV/paiKAS0UB
e7cA+uEw+ksjknbV4UmDPLJhsAmBoIUtGEPzTahDgeTnzGRffpa/M+D3rQVC+YSj9NF9WMpjkXxK
w/dE2QQPld47c+9QXPq+4mr88NWi/Pk2WDLvaf3PhwukHEhASC7kLvTiy0+EozydIwvJ8zD6pmNu
pQIcYlV0CwFpKalFMG8dNh6xt9c4jTF3ZgbMmiLsmhD+TV7yR4aOhaKUyrv4O0c/FfynNwet3gGH
uODsuoxddWbIHhBFvkb/fgl5mxSxgBmF7ARHmfu0dZifdx2QXejCUtv8wlsw0MSTRIAqQaVOlCKf
ChPhni7fToeoEBbO/vC1FoOGwosSb662pbdV4GTlIuRWu/G/Jj/gcFeYwKU02zbQRsuWK93AtWwp
Hkpm33M2b89bXWBjISJW5Y30o3n3wr7sez+AWtDLdmetin1RIPaBM7ULjztYep9DewqQYnwEufPL
uHN54GPCsGweHHLlbIE0fINxOZU7lewrdzhWcrAUl4Rofu8BNM+F0MYUfxPqOz3nRJiDjCeDt4R5
fAYNCMwi1vML2x8zqaoO1zQOeyyQNxgqkzUA3JLP8Qvwy5GNUlhkmRTyEagGjMXcXkzHQ9zNg7Gc
rw4RUg/v9MWAEJQXdvwPZTsPfACWbjc7s8njOnBI9ID6NhcW9P64h11GN7DxSru7plcn22SK41eD
YH4frcJsxGf2mHT3SnDkSHkCJ2VrKlXwq1hHFCh9lMho9F1GT/4x06SGRNGOuOyoM7O1RcChGab+
zzA5pV0E26Ceud7ur9mnDHg9pv7kk9uVy5dRcCQv2xGny+DpICzmNGv0ILN07WzHr8EPM+4tmqEM
iHySPcm7U7h8GQw4L1lCqX1Cgw4OWWYgQhbkrhJXlXsRJkKdA7LbzAmb6XZ7nf++Y82PVUAw942w
Ozw8hvQQZmAMmie15pXdMRk/8fBG08Z27DAN6jkAYMYK8znET8zf1xGpfWy3hl/5+jBV/bt1rANe
CQl778yDGbOU3pqx3cZoSMRxRQKqyXpdYVrseSn52BXxqJUI3ELJ2lIOZmqclDGdKeLEzDAP2XpW
QY1h7z2asPKVSQUVNKrKpN592ws0zbPeRkEyVUxbuwg8UG2h9SvKDm1yBx+c8LvHGF86hg/TMoku
Ll3uU1tPZvEIL4IfFwVwSXwG5MhaAAXenB60xSn+Li6phFJ5oM5tNWu7dhSABmJU/2XJFO5Dt80K
Fg5e+T/3Op/SRNjIUNP16upowB6z7vFaWzXRcpnJ17Z4/wf5vDbCICRRNA+L3MBNbyupAJELQ2Ju
q0iWd/xfH8bbMSVbErKHqGOClUEni4GPuu1Evlv8Ipx60VIKuplX35jZRLJC+0EU5KPIg1z1dNdu
1Oh9xSALWYkNzGp67F1JE9K7ZJH0SyLNpXK7VLT/cyFzbl2I4WRFieX2UGajr1Ti9oOE+pWxAvx1
kWV3ZHmMBfNhsl1GOD4QEBuVDeqcYax6ZTNu21JJrCp55iYe5SCIEwRkoRwYcqnx1v06+cq5TZL8
Y4AaDvOBu37xg8vfnlVhViEaEBiWlylt/vlJD9cvg9gonQqiA+erzx/VQSD/xS5V1y4Gzn1TDYST
M8urf90DTTzITxhBrp/AD/ElX/huDbdCFqDTZAm7lsJVmKNV2ueJh9VqvR0JDeNvogdsbWEp9A4U
1Bfo5cgMd9hQB/9gQY94OqVXDf2J6p9PRNK+U1U/2R8tL7wYaYpsljuoPowtRh7vEYWOeUv1vlaQ
39rUENXhUKGRdTFGErEmgl0/zNxjVNyjrjOkm6Vb+koC1VgGiA0xSnDKjomncD5BCU/RHxk0V0qe
Oc770k8FxA5sIGwZZurHFmDj9gmKejgwm/e06wECPNbGIjSb1Yxro8GShpDbiCUfyJqp9kep5byw
vMtPad2RdRo28K/IK4uY4BshBiMCwBS8oV3DJ2FSPtI+tB7o6BT1NvdresLAGnvw8cv/BGiryp/V
GUDRHCOe0oPyJviYXRaK1xKTJfroKQjp2vffyGe2WEYrIl3ScUyU7tpZs506xjJB3NAg0uM8Q8U7
eLJNwsvS6PpE52glJdZ89uu4T8reRYqeW8Kn1pgSX1WR5drjmF781sNye9ECVF0V3ZQLdJx+CnjC
H3ANs35JQfK6oP/Ak5SY5IofmO3z7daIp5oysz5cx95DxwCIWpjurTMb5azguXR1rn5BAyJ0Mhyc
9T89xdRYFNAw6UHc6Qryf2RySx23YjdjY26ndTm9KOwNVGUjqG+DewRzZyFGsN2E7a/ou5RtRiu5
CE2kizV7kuZJR2ONJOMOwsvuTYuYTNAIJPOG9yEY1Bu5pIlUUIJgac+A1z6HVOXUnv3LEYX32Ovi
4NQnQceLH/2QgUTenMDUaFDywSHcgFQAXAHPGOfzB6yN1cgNYtmJJ2pC3gWZp9JANo+WBbSFevLp
0d6/pX5GeO4RpsJVlJw7EV1NS+Y6M1GNLlDowt+Zqw2BBaIdu6acC66I4OofjjzlsbPp7xi95TNY
VQjaZfZqrctETsWko1lah+h2S+G03SmlHjSCN/6Z3S7JE4PEofwslwPB+JkrQZLxj2sYdG20TADs
ErRMnrbhJJnhIUOfxtkKYWrS85k2RZcTvSKSz6dTU52XdxQwxmE6sBN/SWTyAiNbcpfaCJvlwSb5
hzSDQnFNwqvCz6mBJl+EzIXjYG1neJG92f224ngNQEikiU2voXnPXm9j+JfmtL39D6mHsr9ueb0I
W3YOcfjmRRDseU9J146L0pVPippANUJyzouEGsM/VWls0sWWKDcfFcHO9ZDeZebNAFbuz3d7zqd9
a/nK26bv/B8J4vC+rsqtdPvMhT+FD2G+fVJg5ZV5+PWZoGW6YzxBLMD/MVRMIQHvs5eUbIIg3stn
2hM3Bmk9cIUwP4ilqjOqtZDytYXZbrUCgviZk9XsCyOSj6/vpBRou7fpTwuQrNq6M/cquFNx+Oxx
rL8ws7DF7YdKZ0g3UNr42LK6VD9fX7W8fqvWrjA/SkbvUUAlURlYg//CjwpiN1UrliM5JFLMaEcK
mtASmMbh3N4JChsNSmbnWgnKjRanFMWnR0hTvg0Wv2t5JSUSuIKlDdL21b7CQYJrdjsJ3jgkDZsu
zDybGCg09P/8t0wAppjZx6I0M79RsHDzzpum88c7e3Iq4m9JX+LvcAExj2OM+mfTqbqclb0cexIu
yuufrs1SZMiOwdKXFl3CR1nr10oV72SntONaxd0hQvMzUw2ny7w71o+a6fkEGpoQ6Pwyy4kTxKJ5
1P5XYC9oGMjOqoe8UnsR2j4othd9A9OZe3OIqLzuQtXNxslIpzMFPkXwUNfCMADKuKh34NzKreNs
04HZzuIEfpwaZcPL9/CfgZMc5vg5SZBzvkcH3/zC+dXjqOk8c8klTkYm4vt1Gud0gJfZiKZ8Dodo
bk1UZMJrGikgRvthqQV61oeSlOLGFmYBZ+3UwTQElcmZxDtyyy69t5LGVhCOCksGIkADqq6XED6J
lwHrPlqi8LTr92tnSAEJUMUAOTFSx/vmjdm8uEhikWxcmNond7DDs8MVN6Yd7DiAu9NOvSPCjJbg
WVxP9Qj69uA6maFwLqIB3v4V3rW/aLE+rM/dtYuZ0hwrHtEQbscHfp1YznEc8qr5u4ARjczEE+v5
o2SxHucpxnSMh3C3U8glwGTtNUu2XMKvq1L54cJUbUeivjhdHLHkJtKtuRiHVNyjoNXtN13XRJQI
vLP3xIAwWh3My6TrYlrGRCLnNh4w0oTi5hUzLIW5sfZC4rTvehTO0SQ9MnFBNQsN87GKGzDDx6Qo
Sfv2iJK/oQQPy8vnqVhSzve0+Y9qAoWNaC8Xi4T0eG6IlaQEPavluaiXlhE+xVPo7J8U5U+kQOUZ
KNMN5vESzSonAIyhEni8Gu+Y+uJ8O4hkwLfaIbLZaWAJy4wdaA/SMHowxbvtqlm1iCuJA76Tpnsz
9FXjk9Ya2YZcHDzGyiwdUePgY6eIt2tOIKbNU2St9ekkorM/u3SOa4lF4Py2JnYH7/oZfLnF77P9
1h/UNbkPzrEznFZ7+xtaawffYrZh7rlL1lf1UdmNb2wfAxKbvSuMU/iKiyC9+Zf7zibXY4Q4rSlj
UqFirDZwYRTNaf4YHBJGcvCu9wvaCe6IzJ+ad6UwyfqqxS3qzSNKiQVWjt7BAQeAfSCyPhoc1AqD
cwu1fTYawDqsAUUm/72+rynurKG2Y23T7QYfy3j/9P5jXxDZKl4LtTgEUYEVLgSmOGQ7tJPBGKdv
B+3rSN8x6hDUUYWz2OQi8SrKliXPpvIBdrNRvabvi/p1G1XAct0wXvBN564cbFyZ5Q6h/ly/tHkD
r7HTFVSGC35yPti9rRcSM7VZVFvscff2P35ac10KfifzlihUTaP/gjB5+kRGi8i3Rinid21yO0qE
ZKhmeSN3rg9jPWsngdv9YU3qa93sROcXuhNKtrebcD4efqPyF2l1B9j0iD5f0jJ1aEiBjIsUpguu
2BFbDVMbjTHtK/Z2wIHed0J2T20ETASwrZ1MmVD1yV77808CmzwFzsbDcaEguXMfm8R2JX3JVyqQ
hX3iX7WgXTx+U4Y7gQzVJ0Zy30Pv07NBTd+vOPdQwLkENtaK7uS0eFRlXIVfAziHN5W4Pjo4IhIn
py8pAshIBCYssQBZcCLiPJ803Q0fDPfQe6kIAw0t0GiDXA3saliFHJiHEAjYuKXEXOhjJh0xCGY5
i5vf4ZBtacjZIT3IjIvpomIKpzt3xniHyg4D2Wy1mQfS0gvprB8jUuwvF0RErsv1oPQ6qHYXSSsi
feXlUZqBBFWe7wMhmRIjFF1k/n8F54tJZ+GM9TXQPZBCJNX3BpS0auQlO9Ev3edTW6tGLu4DgiYO
6R470wGmHvXQUawFTv+377zEj7GcbT+x0f/OJGOlSfjYwDVTfUkMGu9vZ9ClpH0+BQBfid3ZZpNW
LW8dMNhPyeSCr49LxdX+iGeQTQYse+WfAW/8a7LDfsHBUSF644zWxmRfNLD3hqkerrWP1/PxH0/+
jThrp/yhM7VtQ0jzVkXyRmmFMInI0eJlRpCjXxxj/eCcv2vZAdm3sTbbK215TrwypluSuzwWKJQ5
ECRxutJ7VaevkA5XY/btMHkiooL1crxjjTV1j23dHx+HbGkb4r/LIQOme/vpUXyep3dx08X6ULs/
Kz6cEyo0RBK2Op+qwgm3AEVzec73kwRL3QLtmHhDqai7qUV9fxWG4euAuFi5P7bn3NsgJtA37hy9
m7w1wTnztrV6KIBAC3+Z/SqNzgYg9AGUWp9LqKharIBJOnfCaEJ6p6Sjk44dhQMdJN8Ov6o6yIsU
Iup1x+7xQEHCl4hsztv4uS3CDbVjqnXObkOa3WdpiMeKB9nNPibWDbhBAY/YNyPUh1zfd0EcbXlf
4WKxZFEri7QvXbNIX7nVudVItoOLpqXkEX81Bhzjr9ynOJ2wlRewSlwpu/OAXm5lmrK9mZtq4+aO
VzU2BYlrC7shNm//oGYpo7mFtHpmOF5MDnKsZs1RKRI8nE+YN+Xx4akm42vESuZdkBvdH6/weF6T
b3kwv5NnFjYHZL9Pw5ghgsBG2+MEC0VgnJCf9KSCW6duThrEIudMCtJo+wKg6H/lPZ6xCyGW0o31
EulAJPjDaHGSBS5fZcKBapXY8EZcJWia1O4cZ13eZJOXw77R/H8VwuqcOoBGvOEA7Oir269NTaX7
z6tYYVOv+Gct1FuFfeN+g4Ht9Cj8ZObGlE/R1jliW3F1hmc4NMnbapImds1u2p1hNwMePuI0plrK
i23tIQEB0A04ytnebk6y9wXmTVUPmLcaQl6RpNiRPo7iMXBM05QM70RgecmhqnmGehsylefE/WFN
423zDSXZsZiWwT+CCpkDw4L0B1OdYOydOnPAJLl+UNFwxygcP84jUkLoj2ektW48bPJtseXs48U6
pevOIZpjWYDff8ILdvQVggY+Dye8KMn6DHjfEOgZu4m83C2u8TabBwkNu97R56qrwfOHrIk3Qouz
eMrovwOcNii+wX71HkhHx3XNnKKhSRAq1KvbmKUq33m84RWFBode5rVH/JE9ynLF/oTNPbOmYmAc
qxQ8ohdyUb8qBa4er8mGUwGfOa7n4e74oPc1rrmx2LqiWaLbu2hrGXIxgQ3jxFEzw/jC5AoXfyCB
IMRYVgYprbYEIwXcyGY+iBljdMzdBzyLH8zheY47UI91bzvjpAVSwTv14cQUdGx3qZ33r1u1bhYM
xDOBbzWvCBSC9RPdFGg0ct0+rotaJUD+Q4VhyuQUodEEa6fmPirHVPM6oTGBVFVM2BpfiKgn/UY+
7KwR2bV+OqnHtq8qipEPx7OFwCaNTUlRs8LGwbq+UCAzK69/clcu2sqiXqTtQ08X+rf6p1rPplSW
SkD24h09IDqyjfW81q+1EoSNWJQX5c5GO1mwED21QG5vRMVvm/iiVCtGJMd086Rq8Tpo8h+R8jT3
l+kehsA1LFdh0GK+LJOHw4+l0GTH3EDDoKKmQoOKJRtWMo0XsSgC9dDTDRZWdOxCO/V425Q4Ilxg
R3aiLTiQDsz126cEBXbO/XDUhw6LKeEHETgOnW7OR9VfQTC6+bwbjb+aAO6dWm7WacqZDcXPMW40
bd8kTlRFLYVOaP+ulSzt7rocTO9HCqXdfJuBoVhjdoQdamKxYoy54vnO1LXr7OvX5KEBj2jay+V9
r+Lf/YxICFOkmc5UPmh+z5e+hAa7WcOqGsKO+xVP5FylB3deDLfvwouMPnI3aKsSMHmGkqwZ5Y/k
l3MjhMWgPizfbukN0soPWMKQy5AArIZM/fq5Lh+O1xzStVtmwHDHirBEviGmUBhhyHTass1UEJQM
u9YuzQis6SJAlMgy5uT9uBdWbjGUuBsVM/FsT7ZMPKb/ZUxDmvmDXXwYM67G+pYx7w5z66ZpaT7P
O6wchfAO0paoakPtw5mLz8Hry0Ul8/jizDKRk0dIqZ3sG//ExwGqzXWALagAus73y8GoUxqJFd7H
aMV0DFFpgqvb8XYbHFWQxciYZSkrMBR9K7qAmdKPQR2xTOlfdhfGI1qU0CewhCCjM7WYjqGY0pcW
j6shsNsdNMCMWBTE+pZYbkIUawwFRus3qWiq1AbfU7G4yQcO75U0R9SoWkc4AAEoDIAmE/nU8vAu
60jR8dtm3go09QWdyhrbcg4dVlCyaY25ir6mSt38enHlOreAnQ7Ybox5mm1rg9TktVrB6YphGDMn
8wtHqZoatTp5hgfye0rg7jayj3OUhrgBFy3p799zcXk71hyo8LKqRL/dTwj7x9ILqHjuskN/cY/g
lOa9FE//JpluNXzT01fAxEcSrNVDg3zgSraUw08L4U0QxZkntekBjWiknzLvmlCIVTmFHFpNy0tX
pq1HbCx6nQAl83NwzwnsWHwJ3TxziXuBH3Uv1tqtuGulspGf6Zkq+15L6gN1n/x2FLx+LDX+I/fM
sQzw7mLFMQ3Lt8rDwHT6xG9prT2XjCSivVmBhF6hV950hk3NrqSnv2Q+O/27llnXJ43KJiJmYvYV
q94L8g0YCA1HZbCaleLLIzPR1JUaHVbgMWJdrRAeCPH9tS5A1UkamzwDizxAiNyeeqIPTaQF8esf
7FQgaX0+5iQQBljkJMfY3nUDZeYaau8hMxEFd8woO5RD93L9CCVjbOOaQ+cX/EoW3hJTh3WQ0iNA
P2DCLfn/XB1kw4TtKiq0WRheQU9A9jVZi7EsDmZvVP8oBjcRr+M2ggvLFai3w5uxlfl+QTZfTNLC
3nw2uWeVvjGZuPj48AMBdKp+MC9h89V8zi688/7OIJFeZgZ1mqt+dmcf2hTc/GyWrdImu7bzM220
gBTvYhN1KyGae7iqIKA6WgSljVOeppVaFmgYiII4RM4fmdLy/5z1iTgZPkaRjXxa48x309ohSHR3
04a6DizfvhieatA0rNvzDB+77h4U7UKTMf0qjHmH+r1DlrNl+d/7IXt57ybHzxbT+cBGt7jUOKpb
mlK/IfiOxPNcUfMWihHkKWeOUW9rl1HDpT15W7e8HDSFIHW/IGXIpzmUzdgqBjsPxxhYvNRVOIyg
Aup7OR+Ax9RsoIfns9mmE+rgPokFDce+6IuUUu7v5orJjWgGGypAsV70ffyyTa9AnEpEzTD2uKV9
+cgjhMyzy1i8K9a6kT/NBYzgWrBwnMvNh7uf3fyPHEfOoVeobNjjxW9OG8rfhvOw5ya9l88tp+ZY
ReD0FKo0Rvnl3xemT+8qztRsJJTW78bVHd4QlTdWZPvLz6Vek2ntj3vzScU7iYU7L1U2Klq8xR1o
T/n4XqAN/vqKDgN+LDCk80NjNZ5a2Pw1RFi6hMXpjFmSFN8/ypPq+6QcrPGH2hjzlsqcs+0aceDI
GuATB/jeAMcgOpeCGR/7mgf0iRxvbF+fyy1EashX9t7stZi1RQFOWL7xgFRr5W24XDHlGR09SHXF
TqlfYkM66KWXFvhrortgWyBNGjImj6xxfas3coxLnThU60OQ4RP9ekuRMpI5EgRh0wNAML4SYYsN
uY3TJZZSPg50AriJs+F5lsfwwN0XOMwBs+CtzRxtebHsDbexzBV/No5b2FSXziJpcUZ0DTVFW4lF
TTH1i3vpGzLrZ5fUmmQUksrClOmbSuquM67pnf0Uha1sqKipBgyGbh7ytkT8Wc2p0YOAJrHP4vTb
XbOuI24/FDBtV94BT45wYFa9lJ8btDKa5wNVFlWEwAo1Ovmk0fORu+ux/dWVZYZclo88dXZ3Q1YQ
QpubDywA8t4qgskDhyKIlvbTcvNMt5kC0JbOzbm6U2yCcdpnTp3hnk6wFVbgT+3e9xUNMbeFVMQM
R7XEARAzm2CEoPRMKfgh9p/pvNp1oZWiXnwb/gOcVOIxGDf9ug7lZtzD6YJb4BZ6lCQpALl1YZca
mSnPrE+srP2ppJhxTLIhYE1ObqJVIq+Lsagiup7ukFtwxT1thkosOyKs87q5F+l/lPC1O1nuJVtx
UOZKVdI0rEFR0vorMWfIjrO2gANAsMEz0bbtrNh61j4lJHV2um6mYaT5pOV9T4eHTIMQLIaK12w2
egpbF1TVZvDhKtgD69FuJo+QDaL1KvLH7eacdpj3jMr5Vb8RvL0LQrPE2Kg59R6hpoYsWdPk48Yh
sr83xislo2jLx8Ow3vTKpZYE59pGcOFbEOzS/Mao7Op225fctvIQhK7Nkmo4eLlnkfPO427tLv2q
bjCI5FTCJfUydi9VjTtyHPnlGxmLvudSwJwdeS+rQt8E6BzheHbrHTSmzYwr2MyXAKGsw54ClWCa
zzTVVvKRd8C4HdqvK3YwQEZmwI8/TPT6ziD9dBOCcZh35Okn8GKGUaGYrtAuL5k+K+QHSeTtTdbu
8r82j/TTK6bOUAM820P28305dXmAyD71VZwCMncYdOYVo+S/8VViilvxrgcANcn7WpC34jn7zySO
7IYCV1IO5to5VvkLSAeaPl7C8jTId7OYDO5tydYWzQWfbPZfpkz0fTSHt4ntuiPmiuYWa1436FIc
ukkhGPT5WzCKoD0nCprOjUGeo4x/a5ze2bmywxuLjH1UB4BG8Prn0HUvUmGxETzJSzL9gunNFAZ2
YubjAbasRVpy6Lz9CCTOzymqt+sKCNVoHh2I/IV25haziRbaeKDTPsuzDro2LTog0lav7FuPceom
i6AXElPsBJXiaDjP45KLBYKPeaGVmjjmnlpEuoLKqrRLCNZdcy3sAAloBun6/ejYAU0p8+uXV9Yl
+3CJCfTR6v6GliH0eMWM5PYcWL+bh8bSxPSD2bo0N/fbtKL+5LHY7nFNS0Kj0H4+i+xmNcdAFYKg
wj8AR0ON/U2IFlkr40+VOngYKEouga6i6/WYMdMOdNOhNpU9dAdgqjeQVytKbA8z93Ps5LyNhU9e
g17VDB6IurgtllyhiTyGW/ycQ/aUHamhfU3JqFC6GfcIC3xzzQhUphVT7L8jnvbzXrIKoyOCj3nm
m1athrkU434VAKmUKFK5Om3Mrzh+/Ywt8b4sV+YN2KLdHA0z4DxfBw8QPHTyUN3Ko8OQF1wSzZHo
Qt3FM39ACeRpkxYdvNkliKz3KDS6Icc4UOwchR29wrHbb3zneVhGB+CYgFLdIZjTY05QGUgKToSq
pCf3t/kCWYWLKd+7yypt85dK69kRPyS/mkkS6gXd3LGjwsPMr+EHc+iwY3sRE00qk47GCRqvuRjQ
2+WZ6ExGfK2gQru7Xe4NN8EIyO3Fo83x9s0Es6yXUvqEDkEVMWxG5/cTh8qd0lYAAY0xt68ufz09
LD3DjQQyBefvc48oFDTZXaHwV5PSAarCtm88oEyScYrHq8LCwzGzM9RF5xKLsncX02mUDzmyblIR
EjM34eeDDAW9UHzawb6V1s3sqALVUotDEnb7WcY1152q6jKgkXtyGeeKVKTNFSf7WjkoNKFzSReS
cvB73D4FVVVJqs9grELgtlNY1V5zqpSlok0zcr1NwoxPC2J1BRWFA7HeMADa3JbE7VSv7AQogX1u
BPq+7h0AKWxGcOp9OdgV5qyKiIOK8mPWaZxcXwjOC+51ub5EYd3qmV8QHmkvf9hOxOPM4cR/X/aa
zhO9ctiA7pERfRL6IeqtdtnJljbbmJoxUv4Z9nBVr3NLfh1CiWCF65BPArbrpS29NUshAM42Mwvo
esLFxEVakqrj5Rc6sLHiQeFiDgtn6lQsOqM97dHD7/5k7CXKXOJXKVqUnJyZ8Fk/CQHrdDWuFaDI
kxmG6wcVGZPtNYUJF6NEfPOiaXtkbl4VfPmukaZzRpymEcNWZRbhMClkU29Bhb1mbwiCSo4Xq7Lh
4gL7PgrWfrRCfJzcH7tubwN7y6aFL5I4pMrY4vBGjNtUAOl0KVsdAPgVI8LIkX2LkD/DJ7eABFO7
vZyaePCqWoqzC9oeME7nl4XXfOfJydKpp2LY2A1Da1LssbSwqRS8ACfW0MvYgcm1bs99K3gHsCbw
QBfdvm7VlU7hiZ6AL01JqOX8MDLKn79azKQdBIq6/F2jpuDzz5/Biu7V07fTEyFm8JLwaLqBg10z
eEypsebaWJG/smbfziqssMwz+4gDQe3wBPDVosRD2cLbZ8Y1oYL+X4OAqCrepaZByLCjHvnuSlbT
rtE7lCrzIHUlMVG7ehCAYjaz+TrNHxLN1aH9S5jsdLKXiN1F02Dmgl2DezWuS61b3GiUNgAAm+Um
9qSLUzQ7IuQ4SYIJY+2TQzdtgBpQQvmgj8kwhuYunr2Dz/C4g41I44WVoFrezw3pfqT/QNmiEHGh
i4keTpG1NfYjIjCTRza8eqPnwXKET3v4OvEUQvlASACz2Cc72UeWIOiS69WlCm1/o3fvhM/Onw1o
6PYUOzRizX7EhCIyxk118W1n8qs6M2nJ5lAncXqw1p9YCcDNgPquWlpE1zvqh4tHuHfyFEqQBjK+
O5o7HVh3+5LWMsePejbJsEtbsl2HwjaAuGCa8ZWitCQL1n/hXWY5tpcpHN678psTjEFmjs2Mfs8s
VCwXAJLXnF0fWnHvFDfnUajzD5DYgUOKMs69yjVk8vld8/orIhxZySvRNse5TqaEhf/b++hIIVt2
5bzksVp/f165GVky/ZVrJlNs4flzhlzL83sRLD4FKWSc20FS4GLzO6aWoy/BLcNjkwMtE2VmHeu9
dV8bSdQUPxv2Gndhy//CvmrZWe+uZpl07RkjQknKicjYG3tpq9umr/XdhXn5KoSncyC/K82sGWHY
6Io0Mcs6DeAm1GApDh6AdPVHsenEc3eX/9/YTOXKPzNGBFGjpHRcV3YQyfNSppRVHDLcm+bSWm6c
svEb4XINgWyYcWmVOYXWaDlyEAck0HlooRTdYn2oTVYtp/5Tt3Lb1WmltKAMg5Ob6x/MP/gzJnmX
cw1Tdstv0gKby8jHH5UL+JUiBqoo0KL76WF/DjENqQUB6QJ11eYceouDFGdVE13EPggQjyRwJ9yz
fSp2JDPWw0Slykeo472lhWTaKIdoUTIvWKq9t4aH4Pya7Cp2dIg8gw+Z5vvS/KGhxSMRjNBCDhuV
nJXKJbs/PQvQxhtyUxDe70tKXMMrvuQ+HPT4rJp9A6iOPrHZKYIiWSDLZ6IkTVbirbw6iF3uJpBe
qBa6otahdofBFkIwacj2z4xJQqOFkuTXYx603eixl5k9NdtflAp4Iz3vkgSJXH2lPwED0IMoXYOK
nl67d4EzcPY81+J47pxCZ89QJqkHwp0p0ZuEoriXYWTmz3EwXwwIQPxbkweJh1w6UMpUvv0psJps
rPL25MhH5YqwTxir/nPDuTxr4mKq5qILJUxUCcnDTLkyF114G3eY41IpXIOuEsWvzr+Ki9P3wxgt
XhjjBgtHPlHBR+rZKtghkD3jnauIb+sodTP0eiWw2FP3W2nbxk2QAsAx5T33BmzcbqS7S8ui1gTn
qjW7q9kEYDG8F06twhHlG07q9WEu/YAj4YuLdu4Pr3SmGSL5B0PGCBn1y+fHjiU75xBPbaivtAsp
3NYOMXMdzdl9rRIITxyE4DjaeG6dr8DED9hsBMd12/qknr8C+XWOTqiF3W77p61pQSFIxLmsE8HE
ol3lzbGnpAcYxbls4FenV9S4T2NJsohN5NK5NiEMG+rfoXq/wDKkklN8kn4aFDgF1aBDUmsuhF57
FXCCB5+hWMohdftC72ZpuO4QCpX/3YOsGZdtcanbfBCyeUiISsSEGvHxQMxkHXCaAUqWO1rzekyS
yYA+3Unnu8ZivAQ2kdS2Kk1hLrxHNM0oLTk8lFFMmb71SaUBtk4sTcWN+E5xLuqG2kU1umaj0RlP
HagPMRbBZGxfH5e0Ps41jYQKZ1UeFaI3dAuC1+xeoBpBMA68ocOwZ28CzO8yx45zylvYSRhX40N1
ig4i58mgOLjZD1VLVBncbQaW2FGYrvJGi6Fw/NqJMU81zoukUAtJZg80VOuCkS5V86M25vqwLhU0
3QhubcGCKE87F4YGU3ZQyiq1mUWwjxZGqSzV8VroDwoEFdizNP7B0bf4TEwVXP2KwnIS+Se7Toqg
OhsKNx/+pj7s5Q7osQHnQOj4uRpv0BHEaqoPKxjFDAz8iLMKhaIVb2Y6vrsKwlcSu5tlE2bdkShj
dgoAVZSUSqrzNlAqcm0xuuwQo7YyLd7XTmkvgwo4Rg9yakDRnx5nyM8azA2U2sGGj+k8fzeQAIeC
5zt5xX5N98hJZDK894DV9ysbEbBFUFMOb3T4sIM3Dni3UE9HH4yLezbxU0VI4+G0/RMdV5WqAqhD
pdcWV8W9b3J5lfrSFC9c5W7qZLysXg/z1glMf7kVsqr1hUv7wIEGtw51pN3SpqzyBWvGPiCpCdgQ
NIV7ID7WaF8R4GIeXV1tm46fMa8tEDf0W6viQ0wl4D3OLpyzO7IjpMstzO6zfUOeGSOiWvRigG91
yZvQwmSNmzdVRGxKK1SqavMr3K6GyGxQALD/WKuOaZTp0IB2BCIewcm7qJW8daAkP5Oinwg2e+cU
tKlk9nqL2AAgN4GUam3rDGAbKuNNf+YHbgJOHeMvp7RWpuQ6Mq+onp6s/Fs/uroaM7GkuVA6LFTa
1BxSYybFn1ay/HL3FqwpXrn94amIIMDda+lsS38R9w6xNC6g2bqobp656Snv+5H9LtBMeuzSddP0
YcjalkUwzJjvmNpymr0L2V1nzcP6zvEhumoPHHR5bYEw/p1KNUwjdR32ThzhAu/DPvuHLFt3MXBB
oDCYehvzjAgZePf7EY1mpxEI5QWh9yz7PfW3jne/3PywONJQKdw7K7u1nbKIZ+7TkngzIXHGkr9p
DSSLfCMVkWewMGPwyJlxTpXsSLq6y8CMvpbWJ49KOi2WALhBVK4JnaIsKeLXVgX823k4w1FVPkR5
43UHIoXSAHYaCiK5zSUaTvzrY0z+Dja+4rKpxqO0QFqTeFkD/tJ09iyvNOR71BCZWAiOYF2T+fm/
hl/GY89I04624N6wRjmX2cvx31WZIggUw11tA+Y9h2OMaJEqJgDNPOXMX2zZt8TUDBCAqAz6KTF/
hbE/t+/qC6BQPLhsipMji6r6iixIRd4nvK7wrDzi7PZuCPxfOK1XWkMr3mQvKgN5IaCDrI7EPXyA
OKunwGt+iFYIHc87OVNUc54ecJBaSK1eleQteV5lGA3qHRgWZGeVePw94V/3yHAvpZ4IhNH2SBBd
DdX47oa3iASS4M/B6ZJ9IcTBSt61X9dt4mA7L0UVlIMhoH1m+ku4SrxqIUNBmbzQdRrsPwGIAvF4
vSFVHa/lNnThL1KmD3gPok+fAWsCL9BukpnUYSZ7GVBfYi8TUSooclo7W0LeLjikIiUL1D9lhhkP
8i28qn1S3jiEbbCY59osvBHGFSu/rf8AAEJR8TBrZAp2I4hnIQ+r9ZCNduWlyg/HajyX/13ykPL6
RGiNBZRCqspw9A2TliBJWB34xEk6H/k7jVEpTyrIJeChjc1kx7r9BdnZJeB4QES6hpIPbnzWTprx
reGAoklTa6F60lSzzI1uRCc4rQlbsn8DD6bahiIhFhxn8oKZAlbwfHTL1r/0GtoEBVR5V9JAW0Vz
JWOuSWKn8XfUbZtexdjSeDlXwRalLvCKSaMQihD+fxglHaJcWV/FM9hXfRYUXPYNcnv7ILJuPGuu
SCd2CWz3FqA5BTzdaW1WDFvFk4+u3MG6rLVBgYKhIVijJnifRB15dhTyZQTLjEKtRVX7ImL+iGg9
rfSjwkOwm7pl6PX+Kn9qwBxt9mOj7Dy6NUNdZuAWC0Ff3rWoYt/AMx4pVmBbpDWgkQO7GqmkSYhG
dSsWzYWunORZu0o5H+fAtixrR92XrXxMI2nolExZeCaXkxFuMx7KTTsi9XFCINZ6Iwt/YUIT8Jc3
c7MZC434lNSSi3hXhqyWU8IEkSSILP/HT7Eng5Iy31XZHrq7bdViwCm40MO7oVjBzn447KZcY34D
f/CWvdZSAIrmqcL4UPG2+AUyF/ZOoFrMn44dsNEYFPoOS3nzfrEp7BHI0fatdV51JBzUfU71g8X6
CyZfnGgEZRy50WmaU6BYpLqdncAbuY+PxgmVjrC8yrrTy8Pfzn7SS06lmuT4qnlQ1lG4+ckoRrDm
5MIdAcYIf3aqNxpMCY9OZlwDEcqdDI1gsudG23I9QjVluSU6J0fgymeYf9iGrljRKk4t2TbUF3/x
WxHtNW+OKmE6ZUPteGqCYlGYI6o7Bp4kma8nFphW8k0yGodoXdDxN3wP+Tjhq2qNSN5nYdQOOc6r
rn1Ov0CD5pZ/nKwISPYbOuOIeT//wzjOKolGY2hXLeNRqf89mTbp07q16fi8o3UjxdrLdQTuNpPT
Ndhsqsm38WW8TYsi7uEhFQyhJGmeA0DBNXJZQR8UekZAVzMc4BXy654sCVS3cCoBRBdIIFt2Xl4E
LeV8GpPdDYpjruF/cixtmCuliHEoeRDiFGgNd6g731m92H8BiOGIV8djeuoiM6+ugdABLAXibSji
QeDMdATUe66Cr4DHYJgCK2bzH1OpIEH4Ka/mljz1yz1K3dKYtMihYijDPY4H+KpMdSnjHoiSxWPu
JPGkrvlKN0JyKafLyr/8f1BscB0W/3IP0qi4Y5NiTP1qAcD4j+6KLoeNgYkEMChjJOgwNeNS6OKj
Xs27a9EX7tkCifEtH6Q0JyTz1VWaXeL+GI6XOzhafFgTE3Xs/3JYHX67ZfBnhmJ2BEgeHLGKiFVp
q/LILJo0DPMb5DihkQW35LDDj2jP0sEVs7I0O3MTC81gni0xSwoM8Tmi39hHJXakgwTrJHNGnlYT
EbjHnHNzN8SCs844aCsXQPh5Wh3YUUpjcPMqWoAnD/mysTY9AP18v4+aVGK93r34UvkfKcsF5aPo
ttiCsHFNRxHlYwao+gt2Dobp8m7JmUJMT/Or62Mjt8B2rV0kdPUP1f2eWVNasbVJuGexMqSD82uL
Fo177quFJKkbXp3vu5m/XvcrooeDuWqmCyDHLfzHtFxaa49x6cfNXK/rKogLXn3AhB2+fF6akZZd
/WnJ5jHvjlbFTcb5HD0ItRudQt3nDwysJgdcVUxU8PKhFPwRNFKZH9P8SLf3qIFTGxg/wSIQGUZo
ek0mUaSs2nLvnFzBbfjwELKgPLvctFnrTTF6WqlwyrsKfgKGzQG+6PGrb3vdDs9dG9LABCbvatcn
fd0BNr16WzSvTrLHeUiYuQCclMhlRQGbJlKj9bvS6jmIGGG5tAKqR0bL6SGY4dU0EBzRHAbX1SqT
m0suSyX6m1+134iNJAMG4U5EKBZ1ptZabSq2TLZ6gYGX+84xEI85fOM3+KPN4wD7PAodZ7nRzwkN
6AFVDnalp6FMWwb3NfqOkm5jKtfs1NCWIaL3Xo4ht7w49gJzSEyC5adEn6EDZGorbE+2zXMh0fAV
6e08jdYc7/ZdJJlmtZXHwa9AcFK4u4Ng9WUuZm/FEdJMiMMPQNb6A3mU3DF3042w8PWGn6DmL7y4
LsMZMQ3A0M6E6IdfyBwV2y2Xtq9j9sdvq+iVL2M2p9RYf2OKujTQvkSZcEuqH1nvhGWM9L/9yCaF
dUGn3bcI/8VWFJ9qMILXV5+k2JKhWegkA52zN11AEQ7PEWhpC5MsZjCO9sxUgOADT73OQKuM5/+o
o5zX+rq4RueUj7PAL+LhYZZ9dBjw7q3AFnIWAdTkqt5XuRa2BHhpUhPmS0F/dXf8005K6LduOgDr
XPRhmrbXN55GqDmqNj+pnBi0QYa2o+A5bjOFehawrmWMxwJq0zO98CaUPg48MnoHYtDf+m89HlK3
TA4uIx6a5mROjU9ttDPCZbJuF4nQiNjqSLA5nwJfbGMLJQd9DTn6qg95jNHmK7m5Wx6RwY/dlokJ
FfoSCZ+LrcGd7cQnzyA+XBaAYochQMgWoWRf8jdMJd17qCGbeGTFdBKMPwL5rTXS/3e53AYsCyUT
40nVflkc19MncKts/G5qXbRrKZhl2lLHd2Zm33dz0lD1rl8/B4+qgWkPzJEALiJxaaN7pPf2q1qR
FF76smFRVqOIBVeh+0gxHQLJwwsRiD0SmwPtX8hOThyuXAeOcSiKkbAuOxiXs7TXMwNxuR7d2yWt
xtTOa3tLklrDfRadsl0e5/2PtzWNBjqqUtNuid5qbIjFDKcBU4hVv5QVL2ob8CwkybjK3No6SUXV
l+HF/xLfg64IPqwWNAib2tH+GVxun6TKmAbGDlAzfl9QTgrd4sMg+JTxXJoWp2vHLIToekpuX2rO
pPd1FDEXSUuKl0A7sLhjhnQoSW6KsxvD7uADZE6pclqj9qggv/xMWZ+cicSbiON1gfB9NVCVNEjU
1CUyRZJGj7aT1BRURaT26UwP2hIdtNcIERn8IYdrhotpVY5VuqmtfZtDZCrHgbSWHtPqNFJnlOYS
nxTL4VoQlKPkg1uCcH+3Sf/uqZ1lgGgwuLmIKoCwYltS5q3m+fwayfcOncPY0ycVlJRk9i/fgETZ
o8U1AYa0ZGKndAQVIJ2AlP9n62T2+Wcq4B1obq9g8pkXVW/vBBckQx/pXYF+8o2SnFpqsCfLggPQ
0LjXAPjnoagaNEWXd+5RWt8UppMTYGO7dlfDw4zLursyftRADQrw7JypjAhPPT0Aah+psZzIVnSy
N/2pC1X2PI7Gc5+aKMCYQzGXtb18eDr6EojBRHrtvR/i3DQ3153Mz7A0oV9euFtiibsBaJZBYdEh
lxQGRxL57bbNiwe01wraVqBTjT0jYLeJScAeh+NJbFz1NsApWCRcFGwojYQiBBnc5yIbpKqyu17v
VeJ4FKHGmn33nKu4sYTwSmYQGclrX6u0136JdJq1Wt8TePvRE3/WZEXdNlUijGfrtqYOrjwmA/dB
h6yWLPmgESTW+MWKikDGcGcwwwg5AfQ8/ZbdygzcrQwjzSl+N65zdKFohFMwWiiFdwJwFLiTuw0M
c++ffWYE8iVX1UNQmTa0OMRRtLAezJvB58xdkLoPxkB8FsEgf4rDl3x68pfE6MnLd5xAv7JwaRgT
weDYPO+vTBsAWC65aorfpt5h8heJLFGZhSCv8xWHz4hMRKqq6IEeuQe+hyWVtLUqAHIUfpVFhf1y
MSEqEuaY13JD+LJoQ3erJfwsFlxa6DkQp1OEeP9ZZDzyDTRAvAuRl7sw1UGXg1D7xppNis/FLl9e
LNd/CSbjm2LcjXUvdkpsjsIstc+EXMAvcFjHXQ0hGM7UiGM7SiAfRO447ipR1IYkQVYsAUk2Y8Eh
mg8JMMGcfQlgTyJTnnm13iSjiu6TI0GHhhrpg9KRI17EWnvJIy19QIBAP5+oLc9F26RnIbV0DJ+e
l5juitYY3zW36eG5echnBArUhSDjKDRLjkCUC2GUd2Wp+czynA/T1Eb1OahvHOv8mByMKqjMdYcv
5juO5u81xGA7761Yl8HhLV0+HxyGzr6nY1AyFU24Xm6zH78RLEA5wiAhAlvtRnkMjfVpQZVw2LYZ
zUibySqpKe1HrwsCBIPzqL2eR2X7UXHewoDOZJ0gAL9y0JoKO/D1YxGjwvvkZathCBgORrl/k0db
Xflv6EmQUjhdFxCTmQbbX4v131c1BWbnVNSoMHcDlBO7HaOnPHWu/a9o/loLJGW9ALUdRBWs4gJl
DI7c5RYFmZIVRi3s6A9UhHRR7wHpLosIA6x3finJKWOzbdLRQWXOjsFAacQLhhJzMtMTsvJUfaEC
OltOJVZ85as1fU1G1o3TaWY1AGsgwAcMi7dQII1s2+dipQ/AyDrQzydx7g9KlOH+q1Ksivc6aReQ
zSV6m8OnARjNFHLdYeJvE58TB+FzaSGAElw1B9wnxPdM3FyZgNI+eO11Nl5dnNvWxQPIHkUcQfAL
cGomNTp3bLhUxyzQjgXlSgaJMF6i8EZmeAWfCf0CErN3rkU38WEwHXJK6vbRNY6voGRfdYOUkY8r
e1V3zoKGUUtxwgiR13R/AHjdtGhMH1vOPCXxWzUcP6TXskLZtWIotqAVoOArUAng/fuloceF8qHT
jiPISUncpI7TxoxqAQ19O2fVZU6iYUMRJRdruoIG0eEntJA8sTQNqA3/aqmwHUVbMGpEEMQBlka2
x/iLJfxPamAnTLatOD666Zn42YHCCh0wfC8/7aZqSzZdsjPn6qbJ9cjr5A0rvRDBlUbDcb8R6Nqu
fKMJHQRK79RP5GlOocP4VF234/j01Wjvy1p/AHqYq6v0Cnq4QEVl2sTvIXEIUfT701jfl911vZLZ
HLifgYkhp9aY88bQ18oAP+rqyicl+83ZPCh5+auSNMxrjvfLP05K+zTULobtYyA6XfC6ZPFcMywA
Xg/1xSIJkIlc/q4CYapAWC/5ivZ9FHALsP/UnUk483gW436n4lbRYbuJyAVLUylrDZhwwowLkwDO
kmt7TZ4AjEj9YybQ4rupB8VpTTfQq5h44f5Imajt8VTCo0Dbp2jb9EZaJiOxAjyop1vKW4DOXJnO
L6c4lGRVaHIlokdx5Szbuoecabh0KY9RYFu7/G02BuAHb8La/LA2jkZTbnqT4ffDXugqltwB8xGd
5FkpwCxM8D5ZlQwxrzx+477zj2AldxpJWh1d6zKM1JKfi8xyps++JeTIkARxykCJcwdF0ypOh9Uq
ky2qTuynixcyvgZ2f9yl3CXIvyEMDT9Cw44f0Exuxy8S/o/gkGNhi31XGfmvuQu7jbNkCMHuwsQf
WBq2Z7fFHDKMxlPD0WV9upY0NWDlfrYN96QbrW66Vw9ypoY+utBYYaCyr43Dc9yv4MQjAPmFAEKE
EupYwv8607BHpzl7KinooKBC1smq1qDg6UAreHaaBFkOsFunFmi+k3PCvLzPgaglEE8KPExR66P2
ecFMcDSvsWqY7B2DZrRFSIX5HHAdXFUTHp4211bJDltEjynlk1C1AzM2lO7W+iceDD0VJ+6fR8dX
Fu0mOtvUYznOJy67WpzCirAqRPfuAZAzFMCuENLSB7MeQQSfI5DHe0W18NtFzrX6LrpkD2dLdRqW
KZd7YCVZOrmSwYn+FCKRcMyrn+xcr15ssQSSpUaxDi79z6N86+Bta9T6hFpWpS/F6rgF1uJyuT5a
52jpB3nYkhhny2HU4lRw1kxGAVOWzYNUm35fKcuqqPjJV5/1oPvk5Zs+MYLOFtQFo2a341+dY4YE
idx+bgdFHQlpG8eBpI5QxKjeG5xILSeknf8vHP5EKEuk+ENVIO8EL3hCfm61tujfUXRhMwZL3wfh
QnATKZGIVVlhuNN+nq3gJkcLXQv+IBTGc52B2vJSIhUQ74BT6/y6rAoo/Qkgd3LPXGL4XmAV27WW
RiOOvc+z3ZKFFDJZtgTisLG+xDhdsIKZ/8hQ+St8kC6Ju9bZyyOktICMdJBNDJTyY2XMAkjqVPu6
RC0ST8ipoNNvdata0316R3Ehzs67BHAk9bHM16fpjhI8URoJxa7tCyDsTsZAl3FvzRWBo6sA6s84
FrZbJE4tW6ZPBoaYv3dgj59E/uQk/RawrSXtJc15fYOMV6EQakefh56oVfJbZaftNanzbqA3tkwD
ghGyIismMP9lPeWfmia6iY33haUrypAcoI1raRdbMubRbETrgDZbU91PTkPWJmtgoO8m4KO7fzPV
qc+ZIH6A7rVogir7F6YqcfGs02xiaIJVOj8Jr5DBXeRA3BHjQp1wrX1bTSvM+TpHPzYh37b9I3Gu
1JzhRHXgmJJcjYA28bRXrRS8TLlf0aQtXD+CA54qYh9dMprBMtOGq2EHBMrPsRR1s1GKukQpqOfZ
0ZYcZICZqDYKHcfAz8rZ+115r1WBpn/8LC5OHgALALXWBq017A9Z92XBBxERj7OCeOGd8dwFBFjQ
IitZV4M8oI9CTp1li4zE4WJCNxZ2rK9gvnFEoqHCS1C9hX185KRJNZokYZYdSISMW/HYXiwq/Lz4
hQS25phwdQUy1Qbh+Y6/gmSZH3Xjqsbevi4YVs/V9knpP87/b5f/LCGLni9KDgoNC5axLQoIDXFa
YOrOWwxqz7yCyePb7uQ9yuQ9rbCe4ngjzQZDbqzg1+Z6umMU+7/F3fTTU47hr5yl9M79Hg4N/TGN
4vvtP7TAnwBkh7FVOMaT/cTD5pob/yZnLqwQ/4GohNRS5+qLCmgF3dCAoc4T2081PnCtaBLNuWca
CRqFNMIlVM9q0DuFQS0ky9TNlcYjfS7vHVKY51JTGjuCRrKAMmo2uO5hnFiKh+02foyu5fLWCWo+
vZ2c4pNEpvM18vG3rAT5q+GXcXIUNDvTpd7eMzpzKhskSPLg3MWU4ZXv/N2wWzbhmpNMmJXHT8xY
gbDOjvMDsTjjwgvpUlqqPXmeClQjDFUK/01bwJD2OsrnYBx89iVcNGQKZjy5KGSyk8amm2v9B3nW
uxEd3PaDR3R8k3RPdvfA9RrPWfRMNcsqFXaKblmQHpZUApE5/g3/THEQLriQ5JN9stiQ6ozUb6lA
vTSBaDCDCV8l03FNjvAk4hihoO4dlGUljdHzRTGR5zbnoiE4+M8Js3ngtZKMMhX2JmMO2QnJZGls
4GoWaQ2GYn5mtOulDQ8uR4SOFxXiOMZtAa0lu0r1kY040iUX5mD2yYIfA/WHACzxRNoOB0qzI5xv
tS8yBdyuWI6l3cIllrixgJHyChrI4GCqA3Xi3exj1ClX0Df/VIZM0qFZpttSabRsRJ5V47yGyzei
FyqVrQdg9UJOKZ2+Ucveln7n1xiv2g81JpOs3tqF8isx9iXK1isSwLE2ATlEfEwBH4MJ8NDxp5yz
DR4H3oUy0Rem6zPLrMrs+ZZeRpD+Xm0wlQ7M+WjEq7zqJxGALy80Zz1tEEB7Mj/BhNiKFk7rFJ4x
0HZsjAl0L+GXLqQkrugmt48SCFML9FHmGO39Kn79bEDIrC3jxXlXNyktOjsve9j0viT5PwfJLGw6
C37VDUIEfo7sr+s1BRebQU9RnLNmwF5hYmNOASwXdG+anucD2e8z0v6aQO6iY8Xmkkb1E7I9NfTd
vYBsZqq9zFZA+gKqxHgBW063iRgI9j/nWps0Uv4UaoQoBwBj4OG3JNRCtRzSPr0MEDjT2MkVuc9K
BgrrIl5QSMhf/JfQFL4A3wpAjMVcBAwdAkH8lB4Yit+7eEe03xanFoe3xss/APopG+Iu+7Bup26k
8+Hpz1nWsj4SpCPDOI1ivc5FH82g0wa4f/GiNIljQg9GIje1JxTQ48sRzzNIPyQBRDWZDWry/66B
b0TfF5wRyb7IlqKlTCJKbu86D8bIIbJAmpB0yN7WkZOTObTsoqhnKbJgcm04YA5ElHXB59Rp1Ns2
9TRVnGhMF1CLER8154HI2qUvgslWWybyp6mpNsYhjdz+a9lnYAmlP7YPBxvnv5/yrNWZuVrmMtmu
zZ/Bg2gK5K7QQpVBhkcbdNw62LVTYNPKK79Ln6uMJT31kBYutSic8uW1gZsB+XCnvaeil/zX5Rqi
9HfUVOrZbJMFeRVXo0fma+VJRzE7LOkvdFtsORCCM64zdVP4HEa2WxmrUYGPBLHqxEX2on5XtiHX
gaP51Nmf6uUaw6knAxLaqg+TdPwEPJztprwasGpfndF131AgbqGBsSNOJz9iqtAFjL8mRvAtgD5f
3gjPXR21BtFDFSBFzaZ6ufg/5olbQAjWgfgpwUZ8nZY0ths/f08tnVxVk8JG4oS/UvpThmGNbRhl
H/t3a/BkGLE4sfoPhVikLS/Z4lEbnsKP2CFKe+Pza0iL2HGqC8jyRs3NCesCIKY20fPkzRzmly/v
x8sNy3fGM83RKtYUgcasK8Gjp+VTXwwy1RGzAkWUUbnmc3k5N0EhGjHpoVbjuPas3Onnrbfq7HZX
HVnkSDPKDNx7XHmaXxtCM99VBYZbnpbCBQGDAcAASgbpgCFY3hHkQyYxdYx4DnTfPkPS0D8HErIn
04UMnLSIQObUWQzaZxcJ1s+8MSkqCx5vB6s8XzYiSlKLwX8iZPdaepwt1sg4abrbguNoMOR3gQCy
68mUuhuwFVkL/zC8PK/BxhFULnj4gtV6144tMah0c7QT7KXnVtq0a0Y20Ca+vLuGKHX163ILhoHY
yJDRQ/m+n5Xo2vy51OA6nDLWz1iNv8wfFGSD6WIp9nfa8e/lV50SWTveY2f0ha2Wm9hVPFUfEcoh
xMGaogS2loGeWFbFZCYT4ClgQUaewVwp6n1mCEisMrer4NMwsDM8EzMlhoDJhRa/1RLVsH3wXxMT
Ew/74jt7/Ld9mvfBZHxfH9lUmX2h8TbXDyWLeFlNk2MXaYGXE0Mf7+XURrUAh236LY959BFDdAJ4
FntM6CP5Ng01IssM0UtBozW+91rDw1eUtiqLip662FnOIj/R6AIgj58HR+V6b6o7XuyzyTqxqT/Q
bo+H4HtgZVWfdJBJzURMHkMDdeN8dPxU1+VqD4jwriMaEEJFQcAHfuL2RDDDi0hvghy+p2vzMs4L
UI2INzMdYjdo2mXjZkLn9WGJLfbHm2nHZXZoa7eUmJvXulys+KdC7AvAFZU0CmJxxywsjWiAis1k
sILize1+Lx/RxQCJ+KcNYzk0nbgM8lKbYUhoOxEH1MKxDWP7V3LN+CXOcEve0edGTA3xdyiRZEoc
HCg7NhYrXaQJWvbfUyWUR3wszhQ7uDwO8u3f6+D9HrvQAu3H4NtHvUpEdlQlP7GJ4q044Ul6W+at
8gC5Zrerg7boLQFk4QL52vECXSO3hhRYieRg8rGyqwYMHpniqFD0gXkyqgh/+qLeQbbMvzGev/g1
/UFl9GpRuL7+MWPUjYkanI9ptwsoOYm1Ij9rwuAtjRDpRCymB/YNGdJ8nfumW6m7uVDd5D8xpLUe
JDHRYoNFaiCw8AqD8mOJgXllheMmhi0eA+1eEx77XceTQuCz1traq6/+896PPViXPZTe1CbIaFT8
BIamWERx/vUthR377y3lObG5M35M1H+iGgzgC/ebw5XN0gO+qbH/NCpXhuWcWOLmeGNiFy2EPS63
KQxGUTtGz70M/ItZde++5xbmjkrkuFeBKiIAc67bDfO4VLnX99Fsg3seL11VKd6VXqqz2Lzzt+yV
6WXcaSHXTssdDCpBsYUSUmrN90t8frhdJ/ETizGkm13iOgg89uDnA6g5gGQBmxs6efIBXyyIMtjC
SL275y4Z3TYxgRD3vKYuaP6ZTXHAcNkEErFbF0KHiBmrrOsYrEQZDPa0mnqXHiMiQIbVhhS6YJmg
cd49w+lum0CbT00QtQUWnfqVlda7y1A7BkpRtGT0XkqmbcZagPDkcS6v+kslSnv97P2JoBBdr/I6
Dumd8Y2R5ZXxH+0oB44NVqIR6QWjEquW+DzolMxf+v5MJiz7PmlBaPgdH2pbBBzswuIaSoFxGP4x
P1+TKAfDkWmjuk6ra+LLy38CQTJLL9KXWJjEGmwK43+vha2KR0lGb0zjEnJRnrSyovbbdPRBC7zX
jPdcTbxVbmVG5OpKKxUR3HpBhi5tI5TrHDu93frgepwAPw/8H143gfFbFLqSuy9HcZtpZoZyuCeo
50IXel1UoVmaEwWIQkA1K4YdcDwo58vHkklo7PqTlU1GwKtex0DXv16KNMeD/WQyHMTBEExrWoGX
CC6S5Qxo/Ll3njONiq9BN+7M06d+JGchEtYwJPzq5V+eNyoj40qBhTl7F9XzDhw5UrBwj1X4pnQx
Kx7GLQrwlYZyLVpTG+e8OZlntZmtGhfRps35qdhC3cBPeXVRlcD8iKNE4yglamIpWiciYaiDuFWW
f86IivN+QGlhAEfFLlbV1rY1OUeotHcFeHTy/92Z7unmCzg/jSmo+odZ8J6s/osT41wG33XZr6ao
36Oxw6pcQ4omieEc5QpgmKKPDrXmqllxZqpGixQ8QkVI14NL9Th1bL6qvuoLNIRt/2vt/++qWIvx
RPYv6DkEiMGTkf4VySImiBq7VeiCpSttBjLaIc8Qf677KUoenG7/ubhqAZSjeXYa84kU3CFve7DQ
tHe10lB+vr2qUj7geSBMEau7I47J8RB6d+Dn66Nu8xPv0fwyCk+AuywVp6JdW6F4I7ADQvqXSRnj
XfHMFs1Ii7B7Ysa0QtuTLjmv98DhKA09OWelhKdBJSaLxEV2mWZ60pqJmJ/8VXQ+O4M1XyN7gGum
gKA/Nmfk8jEwcncKZSUTKDOuzUjrbWtZfIV/1NSJ03pk8q+ZI7knx/7ZevusjGBS7HJH7WfaNDQ7
zM17pS44Jekl/OCg6DQMVbQZHLSalXSOWTZdUOl/KtGd3zPP8jO4Y7nCMJflbsQbgc0zrEyUFF2b
BNW3uggKheJ+CNIiib2yuBXO93lteb+nrubNymTQheTu1f1oYg1UYn03suenzk9d4G2+mMMQvR9g
D73xH3+ZeMEIpKK5GQh8Sc1JPG68azowusl6poj9yCuCsd7VeHcybju5O2vhMbFT3IaPu5dufYM4
bfPDjSefULMFhbexRoeKNcY9xCnB4K9fPiDxar3LT+vRRMUOzk9HFY3QkeP8pJI910LwvPgHOlRV
WCf0y/QYE4hf3psrfjAzmtlQZpSGhcsvM2GceiTWVnifI49pigTvxKWYIXneQ0euW+UcBy6fI6kJ
ZuunUyLlUuOHAxK6h3pasPTYA7Vq2VVQnOKTopduUoC6tVCj0IvQFQgxzw+cf2ObEz6z0e7zJ8TJ
5LxFDkPFulQn0f+iNlPLOcY/Q9KjZvrtpllNX9NitRLvVV+Z41wOdwFLRxAV/M7b2jHKCeZhfGv/
HVa+RgN65PP3FGoFBUVl+MMY/vJGOCkt0KVCSit9bQrWzuOUaQISIhsetApf30sDMqyRNYbJVPp3
Wr8IcRT3m+shSxkFJ/9qhsC1TX6A+0b+qYDMxkgfu9S+UVfsGPPq6japfGNMxk2/m5H41ZFcoMJN
KggGXT8lFC0RSF9klo7bUCKagoB+ZCxMY0mk9/nTjHvzXeRNu0wTVZX8BOp2eBrDetm1oKrlbkBg
eWYlJFAwGPqWWJNvvfcaHLFW7Xt3Qt8n1vhumMSOlF3Bfn3qrIgBw7sYaLrWMg5f+AkUi6n3xKvI
WBZl97wlClYtWtrz7JO23uiPMUc9ENmslOZyOs4yGihIgw2aRf7yItJZT+T5cr/qgBRdJYZXhf/8
WaPnfv6y5CHsrOXQim3UzY39nW+hdVgCgUZHeh6nvofNtp02whK/JVd3ZVMkZ9onY8WZ281xOfNG
SPnZXh6kLYKra5tdwOjzN5DcKkHzdxCV8ZXoEoZPO58IVrY0l75LPW+doOvOnEBaIIdYtyYveH0w
xLRxTZcfAjqllisCt1P6AxuUwpIGSHc5uSURmMULjgBiWKd9swskhiJqkwrgs621t506+BacTIZg
HBpGtX0BH8/XF/HSvh8EPqV3IAMdvjPSN+LugSavvjipRuXwktne25K3vL853SISOJEvpBOuBTCN
lvUAFgGft8o37d+DewCkIVfHWB3aYm84pHEM+f0njeSP2kcEQBe48vepbGrh/dVjYipKoB92hmr6
p5/XgDVKWA1ZSUQMcX1nTr6aY31fBGk6Yax3yRJEUSeRLALRRvjFN4n3Qe09nddyzLFtfNvEnsVl
bHZ770ISNXYmqOczut0ZOVlKkZg+vDooKmdsx3KeNOe1CGZ33LQ9sYVS18T2oTX8bAeNanAoUgo8
ZqSdvHDRmZe3MFlxB2OHVP/7Fl4v2dlsWtnWO830/ba2QU3yUSqc5eWS1BNOkdP4hRMzKX47Vcg/
uUr9cc16zGTc9enfwtGGQw2yquLDeLBw9VHWns/pWmROJMFFkLRDnitpqCeCQBMBauz6O2SkvWms
8rfdo9wMsb4IAT4fqgwuFkGlrf0U74NORE2XLdr+g9BT7lPmhgx/yISNpab9+x9Z/HeCaXwBPGoA
LK9bgjAnOLk0IDDWWhC3W5Ah+DFuzhMfWZQTU+8xfJ4isxMFaFfbkg8uvL5yDOSbRl9uWY/G5+I4
OGqwVqHNs7RhtiKUe8rrkSVG3ie6+NTxqPuqXNiuCeSUsvxyOapV6d6vbxTp+dgKmhpByXrzqyYo
M7p2sQE7UVU/inoeGLndrrGmUKMjVUGXyTukhfLPxp4sRVUNBYfE7dhHsV1XuIZa76F9PmRM0tDf
ehrA9ogME858VxkVNrLwMPtB+hB/twTaGujiUsLZVH8lMlP2P1QVdDiKIwVEBznmMwVOLPs5BWVq
6FrIEK4mbYO1iZ//olK4buVTbjGiBeUJtoh0LMTfrXlBkav2nC226Yq2r/pQuKhq//bfMGKvZjyY
3SMmJGUVPFsdLH/q481+s1XUoecASrOcplqXqkarU82T2PdPDRrt+A+LrIKF0MWYeAEE3NXQ6Kb3
EA6DIZVRVH017TT1roIVUxRzfseqBbbAodA3jnG/W97IzD7ohOxbhpHfTe3+5uKbuTvzL2+ejDoi
47GjxlHkXh1S3KO5QrYRnbJ/0321++Cn6cdCeBQX1bYuisHsNSQJmQ+dz9DuTDzzpK6rlnXKV+gT
I2G3bZ6q8j2Niu+g4WLbSYzOPINouOSa48wkXU0wGIney+FOfXRb4GtIumwEicUHCeiopaPoWfiw
kxU7UF99nvcmga9vX9yIh9NbPRyrwx0dmcC+NIKqdA0j79bxKUCz5dXI0vLRFHsSEixwf8RcFSyJ
fMOEsHG6NP6VTWi+jKIJGlDWRwJZK/N7rV/YnBwHhw+M9PN0upXs2gpJ/KmEZWhp8vHoh95bfTjG
BO7/N1DfSKTEO+tPhheuTk0k4HF39aTg30Mhgb5zu5sG2IbypP+XaN1hCedpJWWHuF+cS+2u0xwR
3gUOeAewQ/VtQLSgBTIzYKG5vvqF5RSirYVBLdOXlbEA3SEvXlv7ph9adGPOKSmW/Sp+fZXtVPe0
MLsXvKPGZYgwLy5HnwWpyaLQSvEVoUMpaeP5h2h0gw1ebd75L1zmXA9nK8NFyZMnSQx7zsgsOpz+
d4MEIn2cFxaL8iqA/kUioat2hq9WJC0MCZZ5tgZSyHfuG5G9BQDEkc5Vb89lGgnj6ogNgRbHe9jk
R4nI8+Y0ql0+tbuxBGxwa12YKneQeVZ18CGO1600xWzxi5aAHTYW4ViDIC9kDAH3dfjIy8GoA7c1
Q/rpZHGijaO3LPNkmsHKxovjc1k25QOIws6fvM4LXBzMmXX3fG4TPUeZLyFaUuQy7FzuoJigyv8W
GnViGAi5H/RamlNFeSPslx5kVYNg6SwRJoHDptR05+O3xNB0L4XjHgPM4lINcC4otimHIwJwR4eg
VHi2A9YKUP9pnTzD0zHLJW5d5bxkCfT+e3e5y8Ee80f6zuDe5MUkVqtSnKeSsTRgb+c9NTFuqD/P
s7DNnCHODoigQ0J4A5YTAqIJRhQ3CbZKw2g5Fm8YQ7Prvv7OdjxOSPyikSfRvs+T131CxuwHxzYb
5Oz3prLxopOn36umppbY6KgRcAp1nJKnaWT95ibfS5Fe2Q97Gjj5KzMRYFjO9Ks/+AcH9dJWvyc5
HpFW8WgDonzv4tGpCwNFqdsvYNfQCWTkIQ4Z1ARJwRrm3HGo8e6c5NKQ213pQ8TXG2br03D+7E9Z
B6NbHkGhk+ZZD1SeqDiNbuYXAdND6wc99Ct6cxLqO7OrBOWE3FOpRpBLevmlDlypGwnvoG1KoTHh
1BTbu30bWTCR45aken9YcmypeQIvnaDKCRR/PzObZrM0K/AcBeFj/WIxZl3ZaUWswA4ERlI1ZjDB
+vHbllDIP0kVsLBaJrSbN39hfjo7aOMHAxyRAghQhhFLwJ5x6lCGtnSIRJo1qwk9rvWyyH0Ci9DB
BnX/RxLrYeAJAsXaMH9/43DmrXLhNrS4kLeUl16692yz8HvcGkDgKEvd/p7wdOnYu1XsUWRwU5LY
Kig7n2jZfC8qsm8CdvSedRtU8iFimvACcaebb4rCyXCOvcwL/iTcVsSQ1Ia5+2TnBTIWJUidxbOK
KSsTCrT9C35wA0YIH+Sx5E4tAI1NKYAwKAhsgbmjGrgI9JIIIbRTNfJZL2P4CMoZEGBH3qWKbCr+
wCUPuXS6Tm8OyjwHUq3Y+qySW1S/ce+VHk49sPMYjSnCHEOrI4DcDeiMKhP6aVKezw6t31GvfQqW
p49lwcf7iIl5Vsz9CxgYJwcZJYScd2I0Yyk8Tr1jEQj5xwXMCt2RkHgqEpWHyI8uZqRjO1UvJSu6
Q9q2mbN95bmYTZ8mxXtO5RqoSX9jkAGnhJpljSVT++s2GWgECXyoUxMLoKvW/On3yqe/i7p1HlRz
m/Fhc4VKT/I9p6NvAxNbsHuWE2r0BFPgrvY1a4Dxx+cVf21XPD8jw506L5I2sRa4cydPupzaO35w
RO62+SuqGVGRwBHoS47fLTYwsUQdSnOc8YkNfQJYxZttbwybeyvwZEalVQSsFobHHAtQMxc9rSdH
AZNM1YJGBIEeKo8szNZdHMbnuVlW0yVgXecd27I3r4yCVC/gW4QJvIIuinSuwl2FcLdfhnJyD4MH
tK7o0qrW0iFJFabrAhvUWEuqdwadaFCbJbRqqhfivYv/gja3IIrWxOUlzP7s7zOlR7bH5N2/cDkA
ql+e+ZHqscTXKG51PkmynQoi0u6a3qU22jsHoHf3iHjKIUVcpD4Y8MTPqB9I5+XNgqbgyRe73mRh
jhg1rrFmD03KMpIX/p2I26MzIzY4+aDe2AlroPjTqUTB5XLUG3YMeedSomQBR8+slX+qqcY5viQo
T7B28FknegExJYNmCf3MA5L8eBU0xHo9vdC2PoQ61/XiM9f+VnTcRyHr9kCR0mCDAiarjus8nsvA
POpTwPBDweaYjCyoL26oAQOMbV5+nQOlGxO2isMFX2zv1drdoN49jRYZPf/TP8adUeZfQGFTDhWV
ie1c01VGn2u8Ui/hV1r6jA5klQ4g7MGJoCD+Qi7BmerQokJFiw474JWipXTbmFgIByQij34YOcec
f1nTGh8YEMcKZ4znCn4aK7MwjX1uP7ZbhGgzFVPdZJ9HUrHraiB7XofnA4JWKX+7RcVLZSjqLxoN
KTXIHPJpGn6xghmKG1ZzgmaA+PIA2cUZflmb5Pc3YxMUxIAkB1pZ3qTKRnrwzq1E7SnO7D5cVh+d
AXYKvFdRasai7FpknDYMPlhKZzjc48gbzwhRs6z+WYZpeM9O2JRfOLUSdhuAqCV4qzbpxZPIv2OR
IWnTafNEO8I5fUjpSZL3pQ1egHhDxpFW4RNPWzXWFhaaYmpzZa9SDD2RTaMS2LyW2QBthJfjRsFC
F5VPSbd4lTcXmXipbJB/lXAiqibwiCOeQ8pat+DPHK/TMG8ftq/ZfvKTakbuS7/CYi1gJ06RlXoz
lOYPMIePquvBru+H+bozXAdPvhyVbR2YJHcUD8JGtJJrfwoYTi2YLqGDaLPxn9cK65JdeWWXYuv/
SYOQUAE383tOD3hRqxkdWiUw9vBkIFHPdXlb4JoK4pHT8e3c7o0tlkpDm+i3iP71xhQeL1BTmaUe
MgD0iwS8gnh22GBq0/KDn60au3xKwqbvy1TeMQcnxDMIc/6dYldT+h4is+QW3EmeLMhwyzRLDYAa
eM/4E8I3zaUn/XKktQE2Cfno0koom3bAU89u9plV4bmdqMehltZQrhtz5GGdPQ+Ftij99PjWk7xe
E/+PD93QrNZnV+IRVreBF+qVhti6FDGBWZd9SkjHl0OdGCjHmiG0KzhSYpt0/QCS0MgELE8fpnsb
nJGwEjUCRu0kL0gV3M6G/3Nc4XHDZ/MdfPcUVtFQJVXN6EYLxF+6o57yEQAAejCdf9ze1foklaVm
3WfJ3x+pjIaSOi5tJ1YwIws31k/zAz6v6qp1moztYV/IfO0zOzC6EoDVYD6htl9OqyJeanRESBne
M36XDntJJ8Sy4zFsAuLZ8vcgPuagBAdKUN0UtBUPvesLiAgh3808+vD8UYMuREIst7S9D+cihS4s
GmMm67YkU6fjmnmoPP4oAtXsJu4jSg/T0ovu2YmDWEy6M+0hO7iVmtray+j/ZOUVYpy3IbHzk9SF
UqYI4180HxTfpD7R/XMpUFko0C6HjTevdvxUbBQp2yJtXJoiEolImsTyeOorjCoBDaPzuSRYQd5z
94cVtPBmIla7ZiBekhXrqWWp/xyzxu2MZH6gXEu7vgnSGk9ctIPCdVJGwbLuQ2glGwXy1GtTXOTn
/+LA/6BJtmPLN2dbntZ4ALmSJiwi2RfG7eEyhH2Ju3vpJw0/I1TXMwE+bbO0re6CuuSi7bluz7hs
FhsLWlAbUY4FFDRWroOAZME6gYW7Hrasd2X5mE1jlswNyOlT2FWTDeRqzAi5gDaFK7s1Mg4vwKKm
tYvkW/r5cXvKKqOq+Q6158HA/bjwyyroGO6LwQKqnSgBb6CcW3JwJeYB9n6zOgiDy4zKffcDwjdv
QfoTCpMiL7TMQguapa/N465GjeG2/fMOHG75PX2/g9/O86kj59k2XrJCvaE7aMHjseeziRP3lkuU
BShVh0V0W5HNNMDOGR4m+UV4ev2iu7L7OXDXmE3EchK8ZBrH3OPVfmofcGMSRIS6JMCIRgKwTuS2
R5C4S90R95oqUtCyrH6QBdGM7CxtiUdup1Jrwz7NzotSR/uCddsYQQM0CUeWxw6v/aIRHgcbO78w
IGdKEnY1kv7aIyvOhsokys7Om4wKVagEHj9Q+o2Vpy/D/5Yswk9S4WzmuNw55xbL/OphyhbCD5/c
FO2aBEYbHNWAzFjMRXX4fL0rEajzlbDaZAmb61JAgz+odns2LaNeVldBlZx27ivfnHVPNKc/tslr
fSTu3mdnbzy0ZhEYT1APNUyYJu3OkmzkOJyje2TQMQZXc/pjpwZ1BzRjLzo3TPr0VWUZzXl8+r11
hHzYJsXubSJsniVulM8NligVIJt6P6E2yknvzyr+DsmAT2u2oi8b7ufcnWeo3S8h+aZK46he7THZ
+OvL9BA3uPOKqJr/lYKBHfhjNwfNhw8+RTb1riTw85Sj2YhjwlrNDlHRUatB6ORRvMGO7AnAJd7w
qWcdspIwktF7A2gfRVetziqFrXlsb26uhqCtKDasvEz2O3jv837MmFarru2MULHnI8EgY4+wNAaM
+XvKvJ0WBYlGSbUnO4oLSmFZe7DiY3XodpOInmuz9znKptfZrXphDVjZuT1SBwGS8hQ0/duxnAbY
t5K8d2y8BOl4rACBTaI2tXsB8/tpZLmMh8rWiEx+X9OBQc/99i520xl3f66jit9Joo/VbHZ15ndi
Fw8j8XMpNH+O8YnZJT5+eF4G/3dUUum//I4t9A68suYtn10et1+BqaVyiF3Mrk7Us5d04MIn18zH
0inpLNFpR8ADoiKNyyE+SpfwtSgppri8JjvhEK5AkEhSxWWU3Zs+84DI11XYpPx95FAMr5XAzjAO
6Id0tt3kayfy4uheIEHV98RxbA8+B4EFzhCHJaJs6lUal4JokcrvtEJWSpFeGB7nIdwhjEDYbyMO
CfK1zAYjmN8MVzkIcwPHNPur+P8K0wGuMDLu/8SILYsqWYaccb3QitVEJi88KPPUQ7ENZ/R4APGN
dDrA/WAwyYqarP7v68mV0PSZzQQq1BwCmElfbg8fZ0x9wbHfI13GaUgnbwrVYJzTG+I0Z+h3VTTj
Knxr/h7aEtqEHHsYHEUumatRmjP3h1yC3lbgxJUddzIziDjoIQH8eTBBjKVXYVIDnlBmiqV4SDmf
nYqcvSgSx344f++H3Z7gtVnYpLVv2BJZITUJDPzpHM84hmPgfUAm7St0CNU7epKdS2MISFec4tUV
GPNN9SqT9qmzow733vfVQNAyudw0qwg3y9S2xCdXJE3aPf1AX8HAt9tjbakfGb4QBLoxcp6EmSQK
iF52gfzmyrWddp9h+SA5v14EIRlFH2t4SeLfVHv6We1XRyM2MEdGdzQvBgnn+FIBzXYeDsogzRqG
srNaWsZ1LTS3IdTvA8vfejTfFYV5WPZiN/s21zy/6FSQ5kwyMebmCoBrYl5FCE5sYLSM4DZEys64
aPtavvpCNHWYdpSXE9PJvDJAj+C2IZegOq3k5CCeFoUHU025/t/i7TWBeYEwNbBcUECW1Atw3cNp
QkdQytDAyX57o1GQfS34h9Epf9dSzZfo88RSHzUvxVaEFFirWD5H246ZWbutbQwwtczttwB3zie2
6DGhNuJ8UIyw8vXOxSXMiakMwISfryNRciE3fL3fkar03MAk1jXtUJ/F1ShLUkpv3ZCuiGO35Sty
kyO7j0Xl61605+0jIPEb6VPtEeeKUpajJeOqYY9aZa/8PH+BmAwFzmALpPrhRn0HpmIpIUuewkD4
IQ4neOTXfpReNjsQfpSlZ5aG8OA7T2ScdYK0kHbw+pxm/G48lTX/XtbcYJvoCu+f64lKAF71hyba
UMOWe7i+xuR7lZKXqoDFu/6PUGFxfFcHYSYQf5N4e0YRCqgz97XhLwv7fcAeg+Zhxs1Wg0HoL/lG
fLPwM26UWNfctku6mMvdMrQ/eNsFCP/r4cw6gGvdAmLuutDObipqxhuqEFkZTFz6TZ1+y8uanWeE
LgsAqAi6YenlTPPrKa8SjGLPfYFvHSslRa0r5yR1HOeZ9pbYRI7NXLdmHm4TPj84RtjJrdWqZVet
swBkaOYWZ2F3INNC7rfCEYVptwPhQoL1Ujk+rBF4suxMVRahk9Afp+oA4cIMN/jMrBXAHkYupncB
6oXd9yyz2CxPI44o3AcA4oxxDCXiJb9aP4KKK4gLnRyJIoOtRVnLh0q2zdjeKNwez4S8PEQcMgrY
UcyQLboPMQZAeXlx0wpkTxbQybytnMirFdxnZUeupagL3qoKv9dYNA1RYEdIH4sKfK4Hz4tlHbF8
pmg0ET7o8+sVvIIV78+pox8ifSotFF7ckvvP7Aeg7IMcG1IO2yXzorIh93gbS0FXtdF0EG96CZ9T
7YriPNwH/IjzWT0KBW8ceayJFzkOk8v0UChPuIPQl4WsbqSa2oyc7ZlICUFZxyrAveFzrUFPIZpc
N43H4PDe6MGLxBvGNFazuWDtm+TIlXdaQUF1mOBmY1S9d5xAFF4pzA9umjdKOZhu9XRLvNvvpCBP
7rqgJDRMkXrlQoP3FnTzqd+oeTmfjXCBYSGPodJKRiB57ZAW8X7t9SqmyWdaDGdskq336Ch/gT3V
5YlOW0wCYJTO7sjFByGzTF7F7kcmOnhUyEdL/X5981bHPb9JZYcQ1jP2fPejBsSTg1uS+RV9IFZ8
o3F5oaWXWVDtjIC/Wf0OhOsI6leFIRniipkphtxblBdoPioO0fo81Kl0zXHwh07joHAOnr0o9v9C
xwpRQYC0zxbmUrZpXNLJecr9sUXIvfYBzZth++CkV48i9QU0DOQvMN/2f02riQpTGbIK/NHHrF0c
2OYoMZ5ea/34EB3jWX3z3O/35gpDcB4DdTNwEVnQ3DWEx0XtDNeswXHVmGrolslEcBNx2ItEBSKc
W8uuxfx6ZbOYkIJWIPNhaFXs4oSp3f3wq+13tX6kzONLnp7lOBuEjsmkCq+vODYK5ekoG6udBcks
7IXQsxLFARvQPQZUly5xNZ41W1xxy55jN3zpPJqVO6uFya/NolAbOA+6VSXEvqrC2fk1ND9TJYbZ
1eQ3es0xew25rrjvReXSGbgHoEZetz1FH1taMtRTeuEnQcaELYyXM7KxhLZY09/r/Jsm7B5VBQgZ
2eJDjWNabalcGYj6iTw2X8MlInoYPTa+Mb/sssjMaF166/9VVxjECXy8RHPMDbaEjuygsO68gQER
k5tGpUDMlPyskH7AiEMbUIOcb5yx6vonzMniiz50Ic9Q+L0otZlelS8yvFcl8HoiBoy66SgRUbwH
sVuFtEQMhs4L+DlU2zbyunyoV3QBM2JODv6gq3DIudQ8fXbspHj+sjarOlaBeZaJ8vGo8r1jtnTz
0M7K60TAZH0lXMtN2QTbF6+9G4S2Ozjgci9FhpC6OCndVsM5/z/OUn7oC8UgqXmZKBFc5Q4e/22A
hvebdcY8h263kW6f6DqdUmsXDd6H65ZKafxEr1liPJppxKd9FKHLqkF0fi5Ayvcp+xc4CGPviP+L
DUjW7cZPyyRM0ywqTUOCAoWLQ0dj7WQz/i9CvPimxdGzGQPhqG5P8OxVYR4wm0/28GFBu/e5OXsD
uYh7zuMxvbBa3SglphxpX9jNlbAocVIVlAWq+Yx/RWaUP9k+/O1jUUnXjBeXSJLbCDRpWgH8oyjq
W689aR0Nkc0K9ZbXmdxDvRUf4tIW+La5LrZX4J5UcGABqDgrP9JBQIHKeM3Q2igcE7yEqJUEN8VI
TwihuHPM06XJWYv8/448L93ott9TWQjVqH/VLrc7eylWFSWb2tRzCFdHKXnKuECfmVTkev0e1iqc
tOViKdopQ87SUbxNPhzTX/ni26NdaDzHKrGrUYuG2teMUaeKnGqFSA2d9NEdh5NktHO0+GM25B/Z
fbJOMtV7+X0Coc7aU1H56JkVbPlpMwg5Nfm/LucaShTuj3wosbmcAPwb3ghxjThsymQT4F2nPppJ
Es0SD1qkle0tSBg8qx7c4fJEJ3T8PXER509CXzL8HyOglbg0NP3wI1c73djhoKe3lBoprf8yO/Uk
jAVrrWbpV4I/wjMhrks/VX2K3gXwV8cNPvlk+a1/fqhGcDM9aP14/okOFHrp/IhhQn/pzUDfmaFj
xGBQIalnGiOw8RnL7CxlIE1hfGobVIctyW/rg1JUuauKci9lKsMG0oKsjBRewxY1aHMYdS2xsTYO
d8twqH9Hc6eozasfmFKr5bs/d8OzH88B4dC+KOdz5GXFGBfkV9lUhQl+TSrNVg4LizTbZnp6eaRW
HSuQyJfoCN9ladmE0ZwL+kouvtTPxb/S4LtHGEb29etey8p8E17HKS8ouDa1gbeweeG64bNNSE6k
2+HtNoV5aVdkOD1oMLrD2KvnngL3Xrfd4O+TMNNdcz72UR4RylXxRLeMRz7cu/UO/jtiKA5zQLtC
KjXYVsI7kq/ih+NinlYLiSyt55lHionbJVq2HMUvngAcFQh64Sx4aAY8kXdFmAOtalNYB9OW+i3g
/53vBzMgZU6N8QA9RWLpT7fL38jd/7pf2KL1fM5aUB4dk2g2qmLFYHGu332UyE9yVkGfi0aIC0ck
1RnjTzgmCvNv7zevN5OovITA8/UfXn3+wGH8tvIknZwtehYO9A1j/36hZHSKkpwPQmgZRQrtCupn
1e1OGllr/UrLuALR6hDOGgTLFb+ABzAeBOaYJYocbcsIB6eBuOOXGi3a7y5pF/NcShDFKojCAYpO
YA6HDbfmejKC3WuMIVTshrA7s/C/wzHdohEP3x75By4FCPysCagYKftqU2C4w/PE0sopaD0v1SBe
TXn2Gwe5Ceq/E9FkgAaCW5l7nLcEPApDyUEq64D4x2V9FZ7hwGOy1yO0En9zMZ28/Vfy+vVuk+Gi
Oprc+wpaMSElPyQIB/TOlUwRFlnT2r0fSNzdVrhup/UHfanuvHU+2nudSYL42qwHKQjOYPt++o1o
kDFiDTbAsoyZemvMShD7XCIn7P4aHVTLKFwUJHt6eqGP0V6l7KKQJkdi0KV6gmpvx4P6gsqcnw2u
Nlunm8rnZpRCvyePK+A1tSfjBPBJQmGLfP40EmcwFi8p/jFS+ISPCWN3EXKqlsf5B2qj0hJUfaN6
wySh55l6zaK2z9zIY1xYBhGZ9ABrGS4K7fDQUaOqypB5xUJjZh0O2BkV2n0d8u5BhKpusOfd4EBB
zsv1q7ZSrkFON8fUpUibAsgEuNbrXP/G9ja8wwVOkJFYxtAq1EjMRsrrfv0rbj4PVzLyHQ4rVXz0
K8pdXS2BFIv7gYSD6Jk4ugi689agbNXErnpNeqPKF93l+oWkqKMdxR8UqD6KANWk+w+D0dYK8ZTl
IUoLfqZy2XNq+bj1lebgc5eLM54vFvA0rIw4G2nY6tLu0PhejhUlmigzwKBObtyq5KuvQki/6YFU
Ig6jS6dugKEYvmqHDfrr7BJ18LndexDAaBWrTpaXzrEGAy6LE4xbyu1lHA+unOpBg6Iz29iLOXLx
36KWDBYhSsh3oC5FSkxnu7vCAGrSIE3MuczhCh4HFtWJduPtpdQiBAtJyGNeNDh08K+utj5D8Lls
GO9LdHvwW1/DWIE8EIgGy923frciLi7T4aRaGx/0SyKpmGB1wdH6A6yGZsVL9ZFzJoS3zoCYB6H/
Glgi4ADgbCc9RmrNEaibCAx0jmqB7cGkEt0dKGicPOjlcOGXTeQ9Cmbh9+PPfkfc/VGLb/JYMX0h
Rx63YJlDhBiNLJ4klftFvMHcDYz9gc+9ksXAuGLnS9H+huFR1TgUBHPN6jG5jTOr8Ridd41xUEMx
aQxGlwWm3FVs2aU61nmJGx3xe+r9N/rkI+ZagACB2/bTTKPoiSYKoty48KpjindMGnSh+6Jr+Juo
p4ll2BrFRztk7u4T2hIPOgHMmxPQ6cZVVeKmcUE8kx+QibJvNwyjoDs0KpWb2wDUO70+Jg232bI9
qLCwHJLwaPqsRBAt/ot1/emAX5nlbIXW0aq+EQpl+96cfBuKSvNR8O6FbQtgDvltqAIop2RxPCrF
KERf/JdLRwVzv4BcA6shmq6qQ0UWGmrAuj8w7NzSG1By849N8vnHmZ9R5Ton/y/QikmKkDutCcc7
vXj5rPUh69SzE0Jwkx200f2ui+mPnALE6dkHJlz9Q92oW1sYsPiOLSWAxW5IkuURde/bLzn8Fv+F
npV2vDYZC03gQUdiuBulhumh39KqdpnCEYLzAaE9n4B+ct2luFK9KiYL9+wAAiyZqVXzdU3iAQhS
0d7hJVFSr1YS28O5EYa69G9E1ADEgx9fyDTHV8APC9S0WOs/NKe4K/xPY9kCZnWkGCSmFU4xgmiJ
CfcCPDooIw0vSecmf7+5Jw6SEnRO38PP0j0KRYr0BHMAgYrtzhpjA16eDCfQFj4pQy3GviZyr6WQ
xI2Nu/fc7lgbgDyB3lD4Y64n53an4/ySJxTFZrsRF0hlVaCIHrQwO4yVfejffRrwKybLoW6nRkVA
oYa/IbJReUf9FZy9O6fQ8jvz4AVlIA7naDFqEUHTwzL6h9b3rs3iahcZ3U3G0uq06gbWRwP51+cK
LyVUEaD87SYhq8K4MNH+KZ3wZ65eP4gjb/Fdv8QjKAal96kc/Gj4YFds7GNlcpu5XmajkM5ran+Q
qWKsgwtAJ5yRujdPcvkAgcAgnyFUiNGUKApGYgmkKP/G6GFZCfrprPUCZYKHu27p1FW7S8XoyQUY
Tm9b2jPQNYZKxmphSKxoPfXYRHtke/uelgMj+Ui7jKFy0nBgqF4lib+t9CpWPmiu3oJcWAQFqpcX
sb7qlTzB8o2NY4MVWqfYlXPZTZcCUATQWC3fS1aUcIyw8cYT+6J2AFydUjZQnzIlJh75vspPHWPG
HwY/BB4PsXRrQJ9S3R9Mff61Cur11t2k7g5DTjQ1G9A5atpl4oQFuHEW7M1Y+4YUx9PqO+m9pBfu
lmT+dEtU4icJAo04ZQZGo7fmNxgBj0MvCyCYauo2h4IWnkVNN/OiFxOx/hh+hXL0DUM/XWfuLOfx
arAcHnvllNw467zJgRj2sCq4BUI45iVl52OsduwLMcJ7xfVXOklw+PPyk4QB5lJVJrP88fZfbTyi
OoYxq8vzryvENhuOUw6Y7i6uy148+fIiwSdshyFETuLY87w8WQFeQ3bu1u+C70hELrcHCDqsLx0C
h+0bYoQKB1a6Jog5KXfy8ubwS6rxaWcUvjF8Pa49u7lEbWBS/0o+JrkeWPMOVdOkLkXMh4SjAEgd
rIv/C8cz0b9gthBHJcm16lA/dJ4owYH9hFX9U0SRgjq06/x9ndXDs/BtjfBn8Z94i8+1h2auJ8x6
7t+iNedHzmHjQYkIn6sLZ35FxbXewAJ+I6I8xFBgoSHMAJ657dINd6DSNFucGG0tPvypeViiSD+n
ch5ko3KSE3KEsxBq9GuES6bChTgs4mD8mv54TQEx2nfd7tgfDv1ffXZRgXGp7gPyv2TjCffESOLb
toVgpkFW58k6jTX77ueLO5ljBCCthZT9nFHB84PW03SldoBOpYdViKC6OOruZTVMx5gFoBd0vKxI
y4iobUsagD4HdKMDoGRWsCd7XvHJ0HuB2IPPbNqbcqxH1WTQNmXaqQhtVz9Pk93gt053VEljzfve
/GF4W0ZrgBF/Rx3UgWu3rlQU+JCk8CIRY0FrYzW7mPCrrwudztuwMoz7D6rSRwawhwP/l3UQHwMf
jbU70+yWAu0XL6pkRgyEUf11nh2gdAIZbgYhJ+lfxPw9+IPTNlGdyelNrrQ0ST8QciP6OzDT8QZk
FicCEHc7Y1jtX5knQ8LpytEssXWX+scIOTlOryDms/z5VCwaJHxPE4cN9w+qEYHtm1U8W+vnFfkB
Gk4wEuGxfhDxunXGUMl4i9MYdnNTFfV2C/i0Jxhyqpf5wmtvPREZ75dNCVzEaLJmLxAJCuF4BIkB
/8nsq26sxcMpHPZuwd6idMJ9zWGcCuZztkzSs9x7Xo1XU+4+GHrplDtrjUzL6gxhdE36ziaV17Ct
p1LxbjDCkk4CwCPZgCAGGlzAN3ZG5HErk+CofMssxKK7FnbMMzqcnjkopFjITk1auqfJhvFXxCfF
CtgzUXc74Ru+CNHm6/LzJkKXmhQpO7KV58DXYLbgP+x7PH5w4CCFmcc5K6ncbfEVSHZpMWwZMvPu
JI+b66nJYhGMJC4aQKWk9joRtPtlSJAkg+k4xQoe22rDRHP8M23eXHQqodz9e+v8CJ7OT/Rp6OPR
UuP5Ht4M+Y14NjfQ2FUZkhGSzi/U5QU/aPBZA2J5LYBzLSu2Av0G1O/CBH1mPL0sEMfps1FUhhK2
vmjfDyLlu2rJVxJG+6pMdGn5v+khpR/MSNfbAZ0MoubYkbegqGyFBttPU90FyZlCmznJKtgddE2R
UbbNasN7HPoBsBHVX6/qYzvLsWqEFCOODoa4zqKbKWhyCKnzQhLT61kIJ5XpbzermZCpbCNbSSPu
/gysYPWES9Ad6g9sr73kTlGMTwsqnnp2JSQrUEgH4w6Tvxnt60AoJBpHdt+TsvhQU5GQXCRkUOl7
G8GZqolpYUTR1Qy5fhKYkTisOdqxlnrJy9TexQ+JonIskeCXI/g2tnE7UJmR6uW5MfgCCT15H7gY
OoIFFzm9ddOlNf/rfYCwbvwaWCxY86yn3WyCkeZwOi6T1gFVV55JDEDfazjuaEJ4tIvvW7oNURYv
rBwvIzssOwkSqusfcCoTZnQ4LaA/j08sGJcXH6nY0yRLxJ/eV3+Xln8fQVQQg7FZUHmp2Hx9LTYi
Vbb5lSyPZ/AYE0wJ0bM4slgP7j+NkzkEMqKj00yi2e4SMG95KaI6pubzvBpV6PVwP7OVJ17NVhTA
Sb9/pNlj4JIp5cZivY87h3NysMzEa8BjASSKGPH2mRdJUGYh5GPKvBsKURYuD5XT3QgaiLEIuaqy
DSK8F4hbU/Vu24PwuLaAANAPGj2blYPjhbCbmTZb60X3ygrPErw4Ne7TJj0bEIl5iCiRUZoWu9Dv
0yycNJ9KYL6A5oMd7VFTfTiAnYxV2SrBM+cPp3ndmdZHfr9JoVtYMDCM6XRJrk8qlqtaqZZoY278
Hd7eus1BBE74MNSCF2tHYEEaNiI7JH2zexDJkafa/929EFMdbmj60WIfPRXUQ1paOy4aVnbYSy5B
/eqXrqZP89w9dl4lwN706iwTHlY6BSPg4mx2eTRWpccmuKudBIqP5dlMXXCvxoatdPpM26F4QSxp
VHPv+2w2ZLiLHrpSsZJKHBkKvzBojk9SG8AJJOJzZiLfSSEFJqkqZ9Dia8x0hQ+14dtAHoPE6qhH
KF1r53FYnnH+M4E5D8k5+vhMsBVHtTEc+ri88yfOR/blaUEfplktQGKhucQQkOlYeXLykfsULGsZ
RbpSYiqYpLvkr8EbUwt5TMbg19NxGxbOUr5CCwQj0VxxqxZi3jvY6/d+YCpyZ0ajqW6Ptt1bqOAi
wofBUZLyusr/akXmWs0fXI78oMeto8peFVquFTiHRTmVL1Lcl3wI0e41ojnQsq3wS5PQhnoSC43D
PUQfeDOVwxH055viPJm/hUU8sFWBsKR7qoG7vgxMClt3Jizs3BCAz5bHSdbpK3S0Q2hGITaDgWhs
q5W+e4goYId4pW3PYwH/aYYkiGt4Ltz0FH9DKzeQ8U5aZcUaLIlztjrVetPuONDPFTKFeikx4qmc
9JEpyVWKScAjW4x5bPGBsEOuwYja1iJwPGYpNv+6k7Ed0B1NkhXIkPy1EtCBYzOb/2fQQBWIMfhu
rGQjqv9V9/blQfJl0umblofN86z6gYhKITq+BXdRbyYCkgVc6UulnQuG39e+7V8ivlcJqoTW+zjF
HGrEKZzjcN6i7WIIQ1Oj4Bsac1dq8G4Be0ZXTk0ierqtaKBDRyMh/8iBNrsjwwaSUxZSy+uQCME7
ZbQIJy3JcuuNGpHg0BZEMtLg8UWQ46LUFduxx+xYjNGiePC2jxbeps7asJ6AaI2GaWXZSJQTPc5l
Nmxp/BGBiSmXWkgRr82yoB+N5eBhFHcPF6MfhmCFuV3ynrVv8GA1Gm95tb23/8ytuS1cwrGlADZa
UXn7n3SCgoO+jzU6yIk7JP+b4PR5JIodWEjosTMzU8uR+EklSKc7ttntLXPNa4K07k6uIphz4dwF
VrTqdzqMNd1yFm9ZdcZUhQb35oSFJrY5ETiqdzJe5Q7zmPIln0cnI7ZLK5Hz6FZ3wesPD/KrhoN+
PNLvK5jxd2Zhx/OxwqPZrGYNm8J9Z0jG6yCFWqwMQQ+wP7B6bKcWsj0wJMCuXTXkS1iEoz8aiEf5
Fl64WvhE6QFZLJ9q7CD/Ay0M3Xbd5aStwKzjx3iGCIQxbAdZuWOQnweCYn1JQ95ZXABIDJnHjfIv
e+rM+Nuh4b+8m6L2IfQvVZl11tA+9sm2VCXFR35rtRCJF7OTEIaH0MFIGC046ydE7SruqHfs0jAp
8BV+7DvooFtEICcbanS6cjkS1Bz0DMboMy4XR+4p5eJYDLgYtjAnj2M2tN6FuWNgEE2o2t2q0Svd
m+k99TiXZ3GYwjCUgcdUQ8R2fK9j+rPB8m8qTWeJLoTYk4Jkc95XPhhYWuvg3n3KUaDe/nFMDXYG
jLz0tEQhQDVPbsglqT3g7W9jxVirOWoYvmElrTnr5Sj4rxAfeAJ2w6H0MPUAqE9eNouz26vOD6Pm
V4FtDPcifFVZNihdLTZujg3UpQ7e8b2K4jnwDR90vCkkQoMjlyVGSntJVHjDb1RvjvIpgXlkcfo2
Ms/qQqzRwRhJQzsUoqUVfy52fp6d3xhaqPWVqJzWwP3uECn8w7wHA4WmQexn84mpowzbc4dfPljF
0aRJaBnTJX5zr1WHGkm94pex5wx6Q8e25GPo4d0O7+DniiZh8A4wOybQtyefmH40Qx0KE4sn8Liv
P4uMI6DRffHDZenOFnLE7SScs1B0azo7h7v80x3WrDsXzL8EbYueED47ixm8I0CL0ac5woeyiXcC
9dZLAtq1Glt4XUeY4H/ghod46QsDjV9HyZNJD3pV3MDcTSfU6Sor1wL23fx6pBSpE/95kWIR3VU6
JUuv4bCCn+DsZNTXIQzq8c4kEKqy8s08U/Y+nsTrzlnxGB3QkV7QmZXxFeAfCT7MCEpbGpxkckpp
jQ7El31xT2atqmvyKTizF2ROdMkhOWiy5swyKBOtFL3Siq1sQCa5V845WgShBTcIqhqYMzDnZxaH
a3UCcLN1fkKiv5XAjy5F3KbV5m7Sa+3vEVmp9WqvGd0tzBLiGO7K7Xzl4dqghmS5puiZuzO+iT4l
/3Qde9Xzpt2AA3VQQCqZG3PNVZtjFLeSyzovhky+EUkUN1dpofs60SQnoGo2gXFqsDlLrkNKQLrJ
CaM/wHY1CErS5Fse7Kzyk8sGHX4+mPEbaNGC5KD/yEkBzqlUZ0BqJlMyQkxOdDD+HD/xs9/uGoSw
pVqLtzUdVuPUgdn2dA2/ktPyVYmCOEYhwd6eQcALe2hUgKPwQro7F9/3C1GRLCGSLqAH7PygHUZ1
CoN5OkJejwNBZb3UnVU4M4klpVFEGyquxCgaZ8ZKY8scLJhMcnWFTHvbOOM9lAAL1gviRUyQBmte
5u0TujoAYrcWA9r2TAqFuzI/dVZHl1vX4YFs6UTyljlCP+TWPJMrUpz2fAoCjgOM0P4BYO4cZtiw
B6su7cpqEz6fzTFfh3605PPP2dFTIf2Qk//iI5AD14xG2gdVGW3ZItx3u31T6Te0Ev5QbXoWP7mu
pYLLZy6GQ80Z+bRmPCYqOFrnJrS8OlDF31kxYWsVmRqPugXnpms4lw6I++3qKGUFdbJqkwsDOiLU
wL+mL7PveQ4glhE9ZzexyO6v5WkmDhvFxFGWHz6mdXFYti6KlwKhiN6KRYeg5cA5piHaNXl4xy9i
hJkBOp3FuMbr8a4yJvWqzIKtU7+MIAg/cUgoNVhvEBGl59FO3oi+5WqMcbJN5ILoljJDoQR6bBux
o9AyISZn3bFgAKvOLWzahevzbxqmK0O+sCZdL7p6nQMb5fXgv7ozCIAunwbhHDoFGT35m71tny5N
4TieoLvu391srw4nbca6l3MQaCqFruYNEhCpb3bnAd0PN/i2iEuek1OVybcclM04AUA2YXl6WUPS
HQc2ZpAPaF5C03Vnv+qlT4l97wmuZwuTuzthbmYSehbPamkCvwBMQC/WO90VTPjUf2YfUlwPXcID
DYGvBSjI5zNn0xcJvTMHIWhy+xPeaZ0EyQ00FKyo2pHRsB7avpf5S1vStmcrTZaLl1UXLoV6D1SM
uhVH7XBPanFueOr/HeZ43z4jF2fIvAUthY8KNbBicbbVuPrpGplLacZ6URHUtqHCcMoUjVIREtTG
k8LknDu3Hrqb+/RMW2o3YjE7CnpkxPgLyijqfgeVG0kTKeDwO0+ne2ihCzgCn1HWMrppz3eLOwVh
FzN5Nx60zgoWPdE4lpbpXhJS3GMBXkBL2M/0xA/BBYj83Th2BCXenPKtbyRwr5Ri6oek9z/Mb+5K
8TJLvdge62oerCziO/C2rN+MkFaHuyR24DkmxAfFfgOr7K5YIXnDuJFP+1dJEXP1ZAYF7I+vSofc
HOmKz9suezuJYJKBaDR8JjKVyfcjrgmhTmnFW24zepvpiuefz1MKA1d/wmr2fQjKBhbzxeS9WX4Y
hjFmWfFIJEcqc49D3S0HFOuPMdBz75BVG0uhI762ExkYLR3+b+y8wdAr8PbYD683YyJim04YIO76
PXkAMt2OHP3X8v6/pAEafj28Rg6cKujNvywuqYtk5ikN3KODD6Y/pvrDlute/HXSCLvuru6I4Wgk
v3D6xxoPIBiAsengmTuDaqSFN0gmNBbiH4TlO4vP+eeBS+Q0y4qS/hhEVJb6aFWLO7xhnd5oeUDa
ULxAsl4x2qT06YE9zB3xi3zUxEPnpI25xJdhDiN/QyoVsR8NuHXYW7rvpyFr9pP3+Zc25Ni/xrh9
PxMRmISLVRXW+ow7u8TX4RZnGodxeM7U3R9IhpvAi5zN6i14eKBhQP2WwxT45/M8OuyYn7uIZJY/
C3iM1sYCEPsDlzkAUvz9zPpfXvsR2gzuvu3IZRIo64VoDr2cS2jUaRZK4N9YGXffDAFs64d6LKhM
4iu0r8tRxv4OR8smPgw6Lx/3ON3mInorI+Or6IkyaE5J1J+ardVK0JBTyHYzZUGqokOfr1NaGx33
yxQIq/J9OSwYIMgftfuZnaIjwazpUp5EX6V20gsACasnpF95cK3yHTeKAB1eeW3oWgmnuEf7XwXV
e4ioA649Aok9/rAVIiQs1NmBu3WRLvTDCqOIfmsmPKahQSoggD4IDgZ+rZHIqXOqk8Cv6KcB+3ll
ozhPDnv4gB5R3BayA4duHFmMs8w+GKIR7jFseHayMqlaSlGTEQWlIDILTu81K56EKRDrWV+14N+0
MrVJb3dl20IcOQLxFzE0Y34/g+mHZL4wa5Fo/EnoCAL3bnzC17+b9PXy32ACM1zVvWuRcKrqrIsG
XcgDOCrdwQUIHND98OGuuPR0V92hzuksAcODYAMBgFthDlOlsQb8wR8pmdKE4C4ioE8bO+VkpPac
e4FM8Prnpaotl3C6LCF+TwEAoKz7QYn6TYSVnjFhGfmD9zog7ayJUupJV952dDNNMxsIJ8su8mBm
aRc8utGcz7N9cwUVjM+1o/NZLm1UdeyzFucAClmBFdeofuZKNVFC9ELxbfq/uIR3PTq8E1rOfUoX
AvHknEfjp8gDj8PYbnWq0do+xl+QfURnOBpHKJPAMLcg+rym23140i5O89YhbgQKFgk5wD78CJwF
fyqOqTbGLTCOSMudPApEwLREX1sd7AY740vMc6piCW92lI1I+vh8rwM8M7GvVnTQSvSzjOmxnZGL
7JJBkpZMGy1EChzYyMUxuAW+UKTCf2tZ8xz50SBZz5CH41sAtLKqTvPIotMNiNyllC0bvw9wy37B
RMNvbrFDLkG7pGDKqcTEnvm2UChGtIEJljIaaEt91dIIWtDUvtMcCBma5GzteOMdmo0gFdJs/gxr
Ci6XBX1oPCWkNvSbx2LjO0pfYDYzoEPgw2LlwDHqkN0H9qn+c1JwkAX31ryPcIS875K3W0c6OQPO
2pPfHBde7+o66lE6SUC+XayUlq5uNuoRL6euKePuJAyMQ4xDksYOuL1OQKAOz7r03J164TUUVhCv
4Cn7OYwzzWHXxZZR7Wwgerb9RjWlQqx6L+ny+pBqrkvz7Tl7p/XbIP/tnt39upMufl0ajcngy3Nx
qEmGox86aBMXbfpfr7jCrxsrtCm/jcT5KHcNlWvU5iDJumwZdCo7h8CHk/ba3mE2oJYg1vxUlulL
ji50GmNVy4WIZSOMo4se+PmCNIO7zPU7KB/Jtj7Dzv5GyTBTyIrEBPItI3E+s1f82bUkRotGGGss
j3G83dALPQrDDlsSMVKpgs6lmksUtesE+cUC6/0W2zWW4Kn21cSAXz5xHQfoKTnDsBzJlnaMUYlB
+BYidCsN/wiG2u2OnuXmMhoeK//YtQOf0Z6gk072xt4TTfcnp1MZQ93DHTx5LgsdWwGuOUE+1ZC1
BiLWXl6YILySekmJnR+SId23ntbo+h62csAYY4z6ZK2CAtOmJbmbezXfvbmi1uvW+2tyqKhDfyG6
w675muLp5h1/qZlu4xYaxCH9ro5ZW6FoaYRAfB1LDbgrQu7KyxTvxmZuXqrGsWnJAVVhSOqmP8Wy
0GaSXXlEAOXRUOTfhnuzRCAoJx+zTenKMY890K9ShYVVLzjX9CdfRqe1PoLE2TptNl87xwRYoS5g
1rPA01kanNuU+AiOlP4gJsQSDnDG4STNCECbrr9Y9lSSNi5a237AWbxgELWaxyAoQBtrbBevx1G5
1zeVQizYBUWWhMGbuyvhvy24H89icA/hbj8fmG5fOq3ZT87sUEU+P3omX+ATOApKn3PW7GYIZVlj
W53Abfrlg97K4CLwT5H3hYvI7qrj035bGsb1YG0m3UoqrOeG8lao5RrRdB1mq0V32Q98aMqxByi8
xSM2hiuMeqqEvAbUOodGdFsNKm9HEQiEBO/XvQXqCm5EnrC1YwLjamUW6VGngu/MnAgj9vhjJ+9j
DclSOr9/EEZtFT52ULqq7RBc0JWG6g0iad9XPHR3HULLeOwbZwKfG9Ccfsc92t3qQF5o7BYd+oLv
0lAjIMLOiQ5K2H6NBLEc4xgkqVf86yVACRzBDYdSBA2KYdxa6WFyOE+g6X1Ovonf5QeOr3Ec8SHi
u6pTMGhSArIYzhk1NXQPJU9hUnR5ppq24WHrQrwcmuAib6zfubuYhrJLlRowasIQvxJzYCvVHfk7
zs9DTUYomEv0QWDXmh4D0nLYi1mK21V9Usbq+d36H4OGrdeiExiJQSUYggSkguskhvtDW7tJ0bYW
X6stGn2kFzAf2P77neq+XAc99S57oA59O7yzza4OtN7pNDozG0YeVWyv4zS6q2j1JktFhEUJpfwO
cixjzJ393ZtHVuJhg03s80BnwU5YtNg+4owVgTy1uZ62qURU4eTvxa2TjNVfaK4/Yq265tBTvMgQ
oFkaftBRFGOwhb6xWQikF93OUGNpJLAGLJ1AHzX6STz+Xemw4iVuzvHVQ7Uf5mS/khnyiJUkVu1T
3iEX99msh8Izlg1L0pu6hp1JLBiPk9lLVEfN06Zl3ci1hfp5Y/Jryi28EfBy1v4fP7TPFq+9GSyy
2MoUdLa4Ny35SxklRjArMnpef0QCNrHljVbbvPU+jsu6TA8Zq86KZziTz95+QGto1VL3h8FSpSyP
819VdaK1n6Hq7ZelO9p6xReR+FESu1WFKp+ssdrxkRTcJxo2pVtoXVOTN25t/TWdfWI+Z3gh8g7F
hivy7VmFSYu18m2LPUpTxrD+F8ChnoEpCn3N7sVTYFd6ybx1h71MaHvhnEluZ3dRd7j8IXa7viJ7
1HdTJW05+3oiPr5HaUwcFMhRcvni7z7ATsFWIR8FLJ2HNfUQ2yv+N03IRv2zrynffdvNzUziylzY
OrF8sxWWYAmBilKzXOLnpCkKlQAzK0rQW+RPBIN3qVPZy0h3Cd7npdGICqQlMrMJmGlb4VY4RTXz
BVBE/y5oKbleVYSP8IbXTEWB7QJ2zc+q+U+az7c1SOMdiI/NgY5a0XgvgJGiKIzt1kskxF9VBVXG
aD2V6NfQHxACuwK++zguaKV+LDvNrIUdHH44LfyD21QZWFsM4/CyGdDyT50US0ckqNQpuoJiYzyG
TNSQTQHFCDjSf+ZeXKFtYWfKAQDk5o3wZFJ4Vf/vgOSBghFirBmtkH9zYLjAmRGmqrwIEVlMc1fS
OoAUKLVOUNyFRZONQ6DS7UOzGQYI/aw8pYJP3QF+fUT7jX9umG6qQ1sFykaWCjCUq53zaiGM8u03
ylM3BKGb6DWbQfSA+NiXFHbFjRclf4+TIdA5ZuztHGbxvAa2WMyBhTW/lgLVH12nW+RuRHsisH27
W6o5H1Ules68wCqlfieeAVUCy1fyWpnoh2DTvUjjaK+6Yu+iPaR98O96bzP9HHCRbm3msMjSqPpA
RnMmcb+RwN5qOZSdQZUOk2Nf3WJiaYfiGZrPsm/DynvXZHS8VMQeGMz/GsIWMGN2mHxQOY5DP+Dp
+Dw9q/v6JxZEm6b3ZXpekUKQ/cq1ZZhWjMYRz+D8CLJFJEavGSQqj0ZzP0iKV7A12JXFzN9w/d8/
HbueQAB7GU7BnSeHG1n8pNbxkew8k3lLSp4VHdn//Vw5JwBTWqwAt0muYFedTkH88jB8xxSgmOKQ
TVqaayLOYFYAjtFGUOcr73PpPKRGaGeWUpbufPWqQv8XHLmB8JBMBJBodLoHTlcVAbJ/Ai5D28ND
xaS1Wmc0yDMseIXZuYOggKOtT+Z03od1tlZn5Y5QVgZpdawGZ4yu2v5hx6XrzwsLWulfFhgOsfjX
fZKwcbJZWYtvBDJklhT32AXot6lyTxuafs5XAbRhEYsLJCPfmAVd+bFXm5W1eOiRbV/yvGEC1rQe
OmicIMjpnPLlLMBcCnjKOtBF8Fmbw/7212xmNNpmndyYfZttfqauAcrk2Mg0ImLpfRvi/AElb8uX
ZdDunZMlyL4IjyWxsIWTZnnStwYThdMXZozZ2dbcMoSUtqP7wdItQPHWubCnFPc9SJxjTKpKsbLs
j7lnDPVGidg9YqZAeI1nTasUPH3Ph2cieEZd2tdsGgB7IDuLfV8ihDIyDL+aIL8JqN5tcr+HnSRE
9rsi8X0TUUWe1ckLlOhhhiV5CzFeU8ohhCSKxwzJ2iRhHCXduyJhxlAa5bh4Dr4Al2xvAR/rlyM0
1NOVPGWgXclJHtlSAg8AKcEQ7/IVQn9W1bkytCaD+NBxizLBiEZPpi8dKz2h5HEYBVck/b0dHMxV
dgNCxJMe8IPPi0lkaqE45wvDf96dH81RD2FnOXagMg/F2tY1AHv6WKoMlUazJVs6Mc7tyXh7V1LH
/NzYyRTJuiL7Y2b3ENgxfwiZHpGWw1KWaNfdjXJJ1058V/zXUtPBLOl/R/A5lHa2z47zoPaVolug
WecheooC+qVFhXAouoNxrVE5L4FGoijlGe5XdDL1QsShfadss7hJI6q0db5AGMM9xvvCrn9Ks4I8
smHnUK7sok836Ni0xowoifDwoi9SS12i87vc9VO4yVyBzgvpGsG2QUrPK5YAXsZFzoeqCK9I71Ec
K7Gj664tasLoROqGMu25yABVW/1m97dt6rivABFd7qAKOU+AH4tcbWisnityA4zaK3k//AVtFlmK
JxiUBHwXEbwBBgfBSZc56G0G8ABGwOppjLNmeR6x4BKrPU/8yceHs0RJCuztQRuTM+PwfiFDbYI1
nTJpSURoJWOKI4awxVYVR9yHVCSavdD5y55YSITHtZr/GPnXC6Pr/My+POx4/p97wOorFooJkS1M
6MXf9DMKVseXfJolqJBPmKfSaCm3kulwZyPSG4PAf7ssP4ooP8pAyEQiw0Kx+TzWTUQ/wr27Tx0y
xLhO+PBP5j+5NJlxOjIh3MUrvl24x0bOfEJApkgvrIws7cQv3psYDXGEXYw5SKFLYjcgGTYoXsfs
AYSeu0ib6Gtqk6+uVyBfZ97hGSpVPRCuevumu1y3gnrOYoC4dYXnrNnNTnujwg64Ok0ELraTGuD6
RNrrVBzgsqMbDHTFE68lYFRpd+VXm1LV/6HMCEDAcVHfu9jJGKou/8rD1uQ+QFEwZTzj/w0jP6kg
9u8VZnEcVFizD7BjR4fosg6Zi2kgXo4yh5GHT1WRXntb6OEEXEQ2W7lC1AeK8wPZ61gj6RokGVwJ
XwcE/5xHnlcYdp2FecXyyFV+D7nbcnXf8t0gLFJPov9BREnW/dMXNKizM1BAFRYOQE7LgyyADco6
os5feapoRiS9WS9xw554MRqArR6UUS16EkZRUvA4UIfKot2iPWWJHwcjjAv9s5SWqq1WQBDAdRjc
TZtj78obmsq4M0oTlCtec7VpAzLAT5zJVsR6UAinibX9GtEdq8DbfIXKQV2ENoqQr3LRufHUrn4N
Kf/DuSul3jFo4ZH7if77mKCd2NCiGvIm6yaLHroK+AtaN7THTgGJnehrQMZwSKkBYL+edPuqtVjq
cZdsocrAr342qsPspModoFyslHoZU5FbC1f4jWx615WfpE5Jd4VO1CiJsyJ31VQp7oZvSmDoo4CD
gtUhvrumzDBTDKsi8hF2PGFP0/Fg2w1TlVCSOQjBE+5HZuoKgIOygwbFxDee/nBM265E3P1hlGCG
f2Uqct0CHJEeL68tF5BhBoWjKu5JPRv8p48o4sabz1Kw4FKNI6ilvy4F3YEu3m0L5r1ZBF6FZQJv
L46c5duQcoWYfndzccc/KVh6/in7kR5+gV1CkLgAx3GwHUNthAKFTaSJGC+v6oOFvnDQyuWn6j7I
Nyhm+uDeNuFTO0Yn3hhRbrc1TH0qkCfiFheY82e9AwfmVJWokMDP0B83928Bxo7k/XTAyJC+ALnx
/3TLqnS2UPvP04R/NYNERxkvW9Xv6ZDx4fuD9qiKKUf7RNWRiljgzdSZxp5YUrgpeqj3Iv7ILTN6
8PHGvazHkBgwJ7YBR8PE0SidR4LTZiqch4QdNE+QYQo+wkAGxxwX00Gf31/7NTh0/9EDQ5S20LOd
yqExSQSnwEcxWGqMOYI4N8xXufFbi+ROaUP/13cnRX6PDSaXMooQIz5l/ebKvmjsL836ZqkA9//1
pTUUcDKtAD6MDhSX6kgwS2BMRr1LI73cBrj7FvCph0dCffK4SqMWCo2+4gy0ws0pu8Y7qhZAb19E
slYIdmw0ICywqwCaQQeN6rMrTIRmimwcS2/ZSzWLDdHg7eKkx2Abb65JOErJjP02qndLVtQR+Dc0
LzvFIRs7J5lcySH4+2t9sL6VWQv/yxEJYrKiJZjjR+hZSmIj/moeoGg0pbh41BmhAohTT9QVuu7v
h7axWgj6gW8Em7bFTCB7l7zZBzpNqKL8csRqdypJs8sdYvuMWxFbo4P472Z06lVneGMrijch4JlB
5gJuw64nPO+MZGW7JUYWMA8bXVxHakKbKhF2E64Nwjk8nCg3ZP7s/BEQlxRG6fwKATFaDt4yyDhT
UWqyor6sUGMkDnXJaiyYISiM2ruG0zDY2W56znc/81PGCdjwcahdI9bZTmQ4Z2b9geQMKFm0BoHU
iBVpukQy2BDTwqZuk60Fsgne6eezExwhNFQME4+YTbBhLb/NEXPqwjfc/tHippH7pNWXJjJUBkXy
C8KDNhlisK2bXDfjRXrXQa1lZtaLom1JMtGP4Okh55nmo2s6fvcYgTyDe0ufuyBfXEp0+9VwPjsr
Cq85ygEF1K5Z4W3CEh2FTp6Hl2/NUgwqjEaFQFIXr0mHOY6D93RyDuDk2qYwGol/74Ov5+X8pfIz
9CarUWLUVw1ew88vGVmKDmgA/TGf9Y1cWxfa9lMFJL53wSKam57J2rsJ0jwyj9evamkSKXwBDRgt
G06kTjx6OsDWdFzJ3uODtyiKDteO++B7oLfnQKuldHv7yUxBlAoauvmoNzSQinpDbDzrl30iv9uy
eeU/0wbrnL24DDm3L469Ax6Ufp0Gj/DGofLhsXB7UizyY5n8IHc5UbQyQtcpFMKNy7IJ/0EiT8jP
eKazZA/EYda5Hv7dpTOew1jPVyIa9npXFj5YJUXC6cMyXT3cGB69kGRCi/DWM3H9QFro47kI66QS
aHIcT0T1X6zAwqOHW3t3R5JP32h7bc6VJBNBT7+onaG3feyStUoDa6I14XQbQv1QLAl4iG0/eLOp
9PgU+JUu20Whzay23RpWiq6jj0etoXxLIGFjq4Q1OezrEKPln+O9A6SlKIyhqzjQ4Ji4T/RjtEiS
bFGkRS6nbdJ6iFfMarl1VNrLy8+e85Jo+n451r2HIsY1U65huMxilc6hJVB11ZvPk7LYfG0PqtSx
GaqBnLv93W3Ob6PiD4MCcQE2fUypgehtwq0vfIarycmtA6Ugrirp2jIGg+TZbNbnuG7pI3RE1WRf
F+hLMq/G1Ksf6F5lko7P+Csmz0XHjoGbvnaUzxr5tGAd7bVBFn4iPddmLLJXaYgheANoXlctxdOH
gvV7dNh2qLitv8V3HOcuoXX/wx6Oi9C5j81KI1Gdv8ViVUeRJoJaxUmO4SUCISLEBf2xadFVpp4S
2XrHuvDRf15Pm8X8bSKe9r3Os5RyZUfGFuc9UfRts0udcfpmLpE9t1f9WmIQy/z9dskPdRy8oSsr
nteCEFHgY/rOs7o1u9NO9w0O+t0ETSuqG7fcvbr8oP4A7/VTCvtwkhNB91XozZn99u3scOiS8Nz8
BfhzBuVAaOWcfMpTFljjsYNFWUKPPnVlj/qho9aI+CGyPE5txVaS2yLOHQ74ZmuodoINPKuv2m46
PfuzfL05vxXciCiLJbeYtUzTaPPtihz9HhtHIvvZQaMHxk/xCkMRJ8bK7vG7D+h6c8LYao/aKB5Y
93z4b4OfxyBOaAJ8Mx06T3nOQrVa9FkNpHd38Le3ElnfPGcieUIjIEHitcVHcVOwmgnxXszM0pO9
zkUNW/K/LhYXNfXTc5DYnncok8xYqYFenfTgfqCmXi+8hRAf5EW9YSZnjxGSmR3N4xUWqpFLYfB7
OelWIzrnZEoGtYs7gGteT9v0uvr+Y+Cz4xI6of9gMj0lEDKUXLCo/R9Jti62YEqL5mJ7OQNJUk9i
49E4bVxmFBAsXEP0jZC9rEPUFFOfxsNfXKioQMwTF4JbDfyo0Uoy9CnE7NxPrqCmt+ao3m4DIUzy
gNhEm5ZSs5YVonLzLpP2eO7RGWZJsHFQsFJLDjBR3k0JpLvqq73CerATc20kAEA9G6sqhaxT8hSx
6GnXaYBg28Uf7+M4WMHR1dczezbnUI0fwKy7oBWxIppu2w7PxE+XOlGEaAJJP08It/OvUSVUWdI7
yJ74NdRbpMkYgEv33nc1qKKQQLZ4wjB93keppBcTet5tZE2KEIlQ9E4h3wTGM8TuTkmk72Lzv10y
cy1sm+n3Wr5zK7VcswxYpWn+8Tv1V76dulOkjlmhKMHQw1wV3Xp2Q+et28Rkz5EJyrFD6xoYyxl5
EHUwzaNS40gshLuws9SusK1aeUPAisAHcFFCO5LkyTsYvJaMPFgV5VKgjazbJ/6CZb88ojeVeYGJ
VyTWniQAhMsJX/XGxqEOQgdyt8BmbTfyMuCN4EeGL9Z/C03fwd5VImTLbagUNyx23i1SkatPN+zl
R/kx2Joeepls0XW4cr8xUDpSmdNs/kZBnRUo/DHbWpO/NvLUcH6mp+3G8FASYlvC+HXclDjQlQYE
tUmst9pM8iFpk0zyehbVwWe4XpvVUkt18CXpPufz9fqfw+nLvxC8EglFDDE2Ub4uzUtV8yoTjGsT
TDCvPuf4iNEHQ+m/lQBk0cNuUTqW9gKElRDzuBgrgAgl/n+BHCX2O3O2a9zhMYjvA6+ZEFWpEl5L
ugZepo+aOjahOCGzqF9QxLyCJf7gx4+B98T06qgie3SJw7XV1O5tZAcN2EvWhpxByGclLK9lnFO9
rhcRkLjIef8zQe59nII7gt9zZ7mKN1ty9mjOCUPBpzoAP8L1Btuze27fGQYqP5cGjFyZ43/OKMW+
cEawR3gwKUpk+iJCl6ifj6kINZlqFTd6/8rk6U4N1+I9+gqXGQ/5J8upwk7pRacc4lPgyM+weyA1
RLregwJ6EbLrvOGJhQGaP0WCHbJlAGWGoSaxeXRWyB+CphQLtFrA9lkOksLZHwOcUUuNSBOc+Bz6
JI6rm6On5l2RtOiSQpUNmc0vkMd+2+W4g2I4XlffA0uYtHr+KHfWf5yZsbo+uLHSfHIWGkpTpKfd
EkOmiE0mJHykAGy9Q7kpyl64My6fr4ECTWMZKRbWMh0FiJEPolfNj/qkXfIq6f/d1Re17yOtWIks
LV3gjEXLns1/gncSt7SWutZjtvxUkgk2mmSHxLte5hrH8Bp9dNuMYKJp5McnF6k8JQ92dStWuJY1
8ezhVgfhHe0zevv/u712SJYm/pLo8rE8bF53S8u0a+JGTO8l6dTIdoChyW9btZGDZXeW9zMhBXPo
3BOsT52bBEx+HMx/a/VIpvpJZpqpbg2U03RvG09VKnwa16SZaBthgFYOpe9uP6hBi8uo9zAh/Bpf
6ARM/q+WEh5UlKntF4+LxFGVn00S/NrkGih9nzh/DbUTOiT+zS4Jlmuov9TUrFqasuXLaGbNIJix
rXwy1R74gl17HyghSMl5jGIVYvx7NzEsNytS7kpaaGw7XDcNB6ULf499zOXE3PVhGwev6hMKNNfl
IQHWzRS95xq1Ln5qq7LJyG/kQlUo5QCAqhPJogHH63g7Sn4MrgXAcWn8uOnAE82qrYn4FvQtk71M
E42ydhUAQfG2aRqdsSnCbxAt+hpIeSabGj6b1CMfefaLTnd5Ev1NEUSW8LoUiGOoAmMg4hXA/wte
LdFLZcpRNui3swyiIrwJeCF2nA/0qjlEcQSNX0/h23FnVQLjlm+Ih9+FOD/3ec2B71a1QWQ84JGD
411/pv5cuHZ9ETmHNX+Ns4eIRzpG4psUTWa6XRnlFuEdFDNQ+1Sypdzk7Sct8i3p5IV5WXkdliuk
FcSM4PJsqdOW44ah5PAha7OvCcn44s7sGxyuGhqPPDSUhSfYUaXGFVkAkVwHIKnQ+XcxdGK8sBFB
x6XQPtdZZSsAfHdEzcNXncJUC/C0hd73nS9ux54rL3dEgQUBOaDJbLP0Kq0rZV+deVGXYRk6wCsd
Lu79vmcwbXOhhJ4IfI8bKsQ//u8W4jVZkI/Ad1s8/tyIJNC0xj8jBtAJs7+RT0SfaiRmc0aP8tqO
cOUm/rPqsVOrJhsl0hEU5JGvwzkTZgo6R+yo9Kky90InvzqtIqjwoGzAmWSEMk2cTpbyip5lTOhK
ng9F8+c4FSJeS4BFCu7LijPLbZixhJWn0LaNsYQcS0PDcCVyzGDwFCAJsTwwt1zoSSZMMCdYsXtj
Ac/G8e8qU6oM0fiaNgktNO+x4YtrYBvxyHq9/4wOwtPhMKPUQ5X91qY+WHdqqRjXr70prj9K8Ugq
pIpq0XykGoK8kd6vCo1zyeT0VJ6Sdf+Tmf7Cq3rKpV/I53bvSMh+GUidZaahZ+d+aeR0ur9fj5CZ
jktVgypqXEWcavcThdW7vw6CdYOXLn//p+J916G9zfJfxOE561CHT5s/Vfkhz2HtGR/pu/hDokrC
NX76N7NyasCbOL6SSs8LcRehQyNUGhIgdB7e6W53ZlZXvNs8b7vhHXQ/7xIbfYscuDdn6FhMhQ9b
nRRfXqYWs/pDG7ArBtOcHf8QD6kRtni/rQVNTfwbOCzofqhVRvauiObLcfEX3A66L2+WqSS9fpXr
vJP+Ykovf8FXTPQkjQwYd1ubgBLBLZ7wOHHeYhRFLGQVtEEQBe04Kcu6e2BoAjJid2T6n2b6GWdZ
vaC8wyff8+lx2v7EpR6mu3YccW/4uRJA38Z6AkqubONSQx7zrF/sCNb+4Amjwt+sT1PpyTzmPgc5
epALHHKTJfDZ5/zEBC3rPQRYa9GHlxaX5A8lqoKgY5aPSWZSgds9po4zXvWknfsKmbZ6d27HhLu3
kbD9aLz11XFUPcYZNoy8I73T7xSJy7wV2Tm5iwUr2Y1e2FGSz5YXUmFrGD4B7HkuyJo21QTS09Aw
Vr92UunLVs0663P4nvneUZvTzE5K1t/Sa1kYvQiul7ZMQVIaxxgbTbooZ0zNprZKeZLsi5n9jeMf
ZB2I7m7mMqOfW15XZWmFbRGsE0gPtO2/18XAAU2Xa+oh26G65eBZapxK4XYSzFKFAzg0KMhaOX9q
HjOlV/T+erO/AYJQXAEw8QDb8yS5LbyrW5DfLSGLPJ3RRZmRSdm6mFyVaZz1gthPOcrRBaN1LMpM
woRI5/lb74DXFy2yHEQ07DzC33PTC80GySgmcgvpPHBSRRH7bROCJgMqjyc9Mnyo4lm5JDSqsdXu
MWIaW+bpWPQHEVZEg9wxF1NLuR8zB7v+2YLalbCjH2UmNW6Jg3bHcG5xGoULCCsyBJB8ypzXUaSc
X9H3m5fLhTY6E6nPPXRrLwLo5yBsrY0OxIJvmTZC4XYCtGtG5lR+iFjrY1R9CA2EifbKYT3XGliC
rwGeBTDznBrZ2MXxoEpcubFUY+Rc4mFavk8Y0QQZv7iJGELvhltyEfpocU+V/V+s70JPyVr14EV4
+hnomZRYz61b0+5xQ7qIYDomrJj2kJjlkdu+q7HwJS+XO36BvpLSyvhYEoaXldjUyMh3BrL/6Hjr
uvRJKD/Vn4sV8pFNpc+/OfYHgWHucjVOnNUox+J3BJqliw+l2zQiFTfmZ3A/lMJpKXPb4ZIdvR/m
1hLoEc6YyKP34s/lla2JWwjSDpPisOuWx/f8XLIutbUvCPfbZ7HyIaJdW1fGqp4GhckbULKQ5hIi
WoLhaqezRGA9HYFZejSchvn3IvVHEvsMnBDri2jSdnan1cuT2nC+w4Fc9DRbeKRl7gPYzSYci2Y7
Itk5NYU8zH2foWPyBaCKZmfCco4SOPDwOljblmbug+iHqMweyBiRZ89FCmB9xyPRbGcCenoBoFpv
sPLPWivnruylQwb//A3EhCydneBX7LGMm9MEhkO95Tgl14NSE1iXmP72Usb1JaUzUGq12O9hPz/9
/XaU2Lp2o9+ja5lQ97VD/L3p4Ej+i30CuqUxMhS5z8I6umfMtOPUi3Z7Y/mw1IDvH2JYg1ryuIn1
5MDiJGPZWht9PIQKNZtpV+mt8Ricaky/cm3HSo4cQn3zV184QdK1ldi4hrZyfvf0krXoyFfqM9ox
guqVUCLc0KSJx5lpNINmmj8ZqKYoqU2C+A4/H3EbqAFG0RYhZa37luLMWsTu5ob7Kof5PEGiD5Gd
r1ZwctoXU8EYZpN6kYRv6mW6XJwN5WKL/O8+/iFNoGb0LDn/X4O+ZWMEgIj+/VP4ZjY2UlQJ8yNE
4AOoNlwP+a1uiz6xfdhEICV1RJTwUpKN9qTlyjpDrW+H1JV3JNp+40oe/5IDPbqQlibbKtdIzHa4
ohQbLUdaoohW3OiyeTrb8PeuCt5CFGnvTR7kPdjJYJwSHtLC41/sstUpTJe04Iqy2v7IUlXXgX3a
AVdr25exQDd+2wGjC0GwQaqJQcLwvrzwvNjXzOS34zYdFEOY3xydUR4YAdeY1wmIrxbxOUzH40yn
jQDt1u94NfxPkWGlxEFNW5r43uRq+CLU6ycP+DPCaUbChG2t2Qj1FsuM0TsvPo4sQedE0gYN3z3d
y46IqzUZslVxLgDGTDzOhfTDXBTUfDw2PAv0LSsst1bc0sQ8fC+4ux2fq2Jg7vIwnykmp4h9IXyG
P7oNWrOWHAOTcNad3E7NZlxaMw71lEwRjbcrRJF1fqRhbDcdeRum46YtZHRhMq3u0OljYYKi0VkM
TrPG+3lPUvQ/vm8zMwdPaOQsAv4yISITE4vsa1Ge8cHr/WD4fe8aehypFfsVi3ClPCPrjZYLlQW8
Yov64bauWqBCbkjuq0/cRTdFhZ8Y3Hgqfo7hmUbJSKH0v+Y5xzQzFqx4joq3IiHlnc3cJzaS66Sk
V0l5tERQlVF/Ssn+FAbsgyxQQzrvmor/HJpUEgbUJKwRr2fobR4RI/x5QFxO71ZjnluetiUnsSAi
/E7c1acjrm34P+vKq51uoK5Hyk3lTzXSmapiPe4XAgdOqhqBHYDFVcvzOzRMLXink4oQNpGzGer9
vlgCC0u3qNRoth/2/+3W/if6xdZyUZYWyUjHNmPazJJF8yonYlUbqpBTUyIikY2ohbJh54lNIk05
RZfSa53ZclkesLBV3dQRBCz10nOpbZz9nt8mWhgkcOzAHY/BytWROdAg3XMjxpHW4mgU/NiJuP2D
XsooFg/KD1mbVprTa82nQxiFhBH22Jjo/ooTGkL4cn6ifF8FM2Cmv90ce9i80gOGMeSp27f4CC1+
NoLIQh/Sc7iILI46Y4gS+TwlmYavdnedmSzVBtwvpxG0VRrPnuM2xgcrqLeRzt1dAEiei5uHpZ4H
CQJxLeRE0aTT1Ss8uYQ7YPHeEYz9tovjT+T285C4CxZz2zjaOevyajCppaimN5jkVBQujWaoRiwJ
LGmqbiT+ssOz23OZ3gY/hxfHRA3UN/yuvAjq5dBVPsPqiI8DIk0phY5knAoo1gPQIudYzUhgdOpZ
DSEAvTB+ppIi6DCmb/2KdsZL45CE4N8S5J1XC6speaOpPejKhJJLR7E0Jxg/JFQIONjUEByIBRUO
X6NWL5q1ljXJCXADqcTJ0AKDj3EJfch1BCZH89neKk8E0628LMHQkmyoXhkzZ5ixzAkjWU+Azci6
KdTyS8vPT/PgBAJysWmRR8+BZTm3cKf1lhn4m9ooL5BlUBu5Qnk1UARiBJ19mGLXlAb8WX/DBb75
vuOy1qoJEkuOIFxYvtlF3X56cR+xz0nuVFwXhYncdbM2X4SC8kw3mwhXdWWZHNgs2q85qk4UPTbi
0OdiICQcIRtb4chw0YhxE4zd/L+hrII1o5Y8xlS4XfZQ8dd9bWdyOfPXSh7uK96U+HajlAvi7EJG
ED7xJJ1QPHSiugN/JjezchPjtgSxe4P+VyGSIxG1ajSZiYTI7JeaNn69joRIwze1PoPMajfhDT9L
1Q2d5mwnSh2pccFfpK8RWfhvXkl+rc8WRGTHkSyhyrkjkCcPAGfVT1SJ+2EoMW4g9+GEw0cpuziy
Va1GZhn+IJQyYLQHV5q6SMBqFzsrgMAuB45wHqSj3p7gDlXpXZst/YwO/032v7gcE10VRfeITuVz
8LFFJX+mtTP8KwG0HBwv9GQxZhXVh9EhemhrTobbTaeZV2iwqbNvuoFq6tfigD3TrniBOqsMbvxL
hii0/5PC1l/i8F3m0y6xEizezu0QEmTW/ZUoFS7rxEwMvhbA3YIIfRR6qnw7IGOH9JN8Pypc9eqw
mLx5zl6jumIm65lklphYBL14URAITEQ2qaTxbYUIIwdjIGKvJ0j3uFq18sSXo9iSBQj1RimTjbe3
rPTq1icwIcWPvBSXZ574aOJM/VvY/JcHYdos/aIH9I+QSggaW80jgr0QfWtP9MafXp8/MOIe/Co3
VH0H7nR0A0xcxyIu5g+1txGtpARXt6yLMjezxsKXZgOlQsPwdFsNdhfrFLRp25S2+w7YPtZQ7bZJ
IV+otu4g1fgjthY65tHCy25YtcKkyNHmOx3pzEBkRed/2kDBdehXsYFSuguXtC2nhB3Yyji8w7S0
ghZNd5n+ob5U2NZCKYPYg7ySzH4LXzuev5aEINu+aqjClpwqD5UANm5Bx+5eW+9A8t1i1FJft9xn
yggjJFf9F+/Qmnrba+BrWSDPNbI7ZHcguiDTG1ZWWSDrVNN8D3Go/K9idxTO9BDcNpprfJCnU9aO
DgMVFcb3c14UcjkJnhVEI6aR4o7ar1S4nTbbnJmiPUNeDwBnB9Qas6XbA4WCut+uLjNPO4TQGnRE
QnbbJ450NCjKWOcAXouIT52UTuTZrt96coZZAvh8wnJsW4mvIuqLSP7FBcosOhuA6viURh9S1DLb
pviYKENsItZUYcnGTHMrHSKDGdBrJlog2BWBvDHApuiHA2ng+XgSsyj1XjHoKdDNLtEFLwE+d9DP
mk1QUxXdMUOJ1WKCWNN4YR/7xQMmX/8/Kxi0cigpZ/JyCPijvNaTACiVEWrJSujnzqRQIKFo1mkx
RKa8FznznpSJczImF+PmDk0YDnvCLxo89KKiwk/R4+ZKmgYGSt+1k+5aUfIq5PHCCeQqI3CeHYKO
f4MK48BapNYkMo204T4liYdP3Eb30zfojZI44Y6YVVAj5OtmWz+Bq/V9RFDboA11dWt31pNIuKuX
8sdcdYFz1neENP8yIcqjn7CERO9JTte0cq1nKMknqf9x2vYKJOQ9U2w+4CFdel8B4mDPBr2DEZcb
bCbAIFLVysONjc8ouQy0Z5fN4+CqXMBasaF2lfm9YQR0/LLRl01iUjf50shtEtIc8dPtwVruMX7L
CYVkFfXFHLGPPxQa4IfOSl39PBB6AIjtpHJGuTJToOIIK4SJxARRAf6+kq5liizUYJjOddY8c1e6
tEEDe8ieNCbEbEM55wrHpZe+2WvNcKEa/dnM52ngsPuLOt/AEJs/CuA2Y4njfRoLYyXgRw0GCdwe
voJQzXOJNbgT44Ey07NV/Tl7iHTRb47AsMrPRK7XYsG1XEenGPgaksB4u0ODeVl5H/qBxvuZeKIH
ypm3E8iKPUzBBvYYpeNqiRp236qsnrfcQzqlfAbYdqqCZb5jLRPs2Thu01Tb9nrNCdraxOY11qWR
FXN0bHBgcG873FlwL22y7qekgqcS3ZIpGeR/3QzjXkrR1RPQT/AyUD2LAb/q3gpCekxnFlajGZlQ
gZC4dR+lJ36PJp804EHaKe/GY0em7lGNBJeDOZuWyvXWuT+a6Jf/dus7V9sVfIf2tl+euf8YwlhF
zwW2+i+whyN1s97mQoK1OqxRyG68kslnZgdVlUq/5RpmrZOD9sfnpuTFotgelFgkRRLgth/L4rdG
FEyKnhq01YpL7UD6yr1WN7hY5/ER9cODY/6qdLr30zQlpccrX4LapZNho1HdXGIo9+zcaie9hZDc
mI9DA1FV57/SzhjeUaqhPdUjRZKBvYOvnuQYGqFqGCcD8R1I2aCQrdll9lbHHaUQxKPDbWOBLcoc
lsMVVgTkIFoL7ehJLZoz5zH96WcongQp3IXUwioIMWL0VXBh1k9SazIPW8sccLdRHCkZBbZpzpiC
Cc7fTLC3nJRhWNnbKDodtk9e+LyUgNPWKdbRsoatxftF1cwP/d+//DTHooQ8ezrrxbudCNCSg6A9
eSde6IvgmOcikxP/6wDrXoAt78xqNzRm6htsVISPu3WTdq/Hn6KUcf77S5vflSGAlpzSwmuXJasn
aE6BMIOaGdmnoH5tsbeZeH5pegHUnE6bQZLSJlYFaJqR5savVkoybM8d9DE6GovP3LC4vF/P0vNX
iL5N5lb4dVQehUDnmwfP0gD3FExjlfUL5B6yq3S7F3+i03PfzIdBvusnLBh26TsbjBK/bXcc5/ip
dJUINxadPyteJtHX/zXEYaDAsKJKtDWoAlUfv6Bml/CUUdK7Q1sO7HfYdRkSjMqaBQ6h3VytrMs6
E+IhKSBQVbZcDC73aHruOcPqm3SgqZeIIe2fuZhJdfjWnzHVDqxwjG7yOIDt0hl8Tz6/E4g+7ENL
6laAKCJ24hgSalBOqqIm7hs7g79m7uJjCjbJDSZmTcKBlq8JszSiyn6bcVXXTAWGimqVHFEga4ub
oPMF/zYtGTiRjaX9SetglDRYVeh0j8IE7as0sVbrxlcc3D44hPAmbnmNV+VM/t/Ch0OgZiE6kXR3
x43rhgonAV4DbkVO/MiKOLqfukB0RSuaD9AdLmTLgIZo6xrHE/KWDlo+tYmmHIFTUQ+sd2JpMKq3
6lmuMfD1OZdfsTaIcgM7qJs4dzddCRswwTEqflmmOaofBvxyFSTOSeL4HidMvDmT0GcM+efPqACQ
lAoVGsD62b8bdgo5VsLzp4b1CFj6U1L2CcPXccqtJpK/MJf7sAaClf+gB/wXJcC0+X6nN+lZeBAD
6wOK6BlZlqRJY7R5HptQjCv9YsVIgpRfDzyBjvX/aid+ZrTBZPr9jxb1QFvywMNbjPLaPaJ53dS4
t6KZ24ShElKTv/Siia9W+WCONx1bU4rRNStzqsY/aax77dcczRRKXfym8ogqQdy33zezo1vidmS5
hyy/Hk/yz/gYp7rybMWjWp/JgC/PrbQa5CXmjUEG+srZprwwRnkdi01n+Lf4RnlYGusNfufs5bB8
RtjIVqDlcaHsXE6zrx5bsGBEmUc1V20AobkqV57XhAv8p12eND/di1YfYjz+DBTs9eheoFT//5ca
PbjTE87LKyuhRZmsmGBsq+XpEwW7TlPEqa+703aYE9RPRJIe4hRVV87eBFi6r6H3jWayvoTOgXUW
LUB2eR/G1MUebEiqGxcl6NMuH//FT7KOG724ad+ayNAYOwWCsxpZj4xY6tRiqqIm1K65L+vMUqWf
90D4iw6ZhKeeeLgPC6ousXJLvLt8Nk6lB8+7Hf60xFyqteyPUO1yV675lCjMTe0b1ET8z3zuzcAC
InC4DxwuhVNRG47dAyUGiT/N7oxBBBABUh/dzjT19E4/SXgx7t4okd3wPBCv7/j/9cZgHMsl68RI
6I2a9bAWX4wUEo+erE20H81qrC91BuvdxiZhlJmvgpcngBNBiavcngwavG1qw/ySuYtMHM7yztz7
msidEdyXjXMrclgjFbxM1cOGQsXe5Hzc8vjWp1WnVgdhM5QbWizH6bmGQ8YH7xUy4lzMzVTJkH8I
7cPKLOwyYtOMAROtFPS2z0OD7gl6fYwoVnC0N3e5Sc6cPiV4eDsnao5VcT1QEwJH8aZmg4n5EYDZ
F0ExJ64C9pQ5rBX+DJwuAPjgQFDnZz9zoNzApfuGoG3dFe0Hyj/XDdKLFklpxzpeCJAmhBG6AeIK
wttaIFvJoNAxnF163NB1C5hYIa5m1hTelFNDm3OHKOO1/LtPS/yHn0KgZBL0EuP5HbXaCwI7dvxl
iGGFLm4Q41Sh6S6qhSBbBD9nC3/NQWEWoSr88SGZQKOeLTw0VQ1CUvYYAyQsCqOtQaVTe7kxdazk
vtRpTJhm2+65mNip6a733qKDl4iyQCZEEW9fCEHSGiygHw0yLBDIC9q/IUNP4EoTopV9UYTOdSKm
tzyZIdglDjtJkj+6uenVjMCwuXl6BDLMyaB+HEZqWE8EZvoZAgnlqpxYVpFopLntVPZsTTA0O0c0
Svd6voOzGI94Ac0bkADT7Bnj5fduOTmN+jkZROyLnBoTgbwjIsBsy7GdRZyGESrdsiRAWHUGHknp
9dPL2ocQYC65cyxEhGpQm5CumuLK+kUJHxF3RLM5+S+wQL4Spsf20nQstStuzTu2mWuvck8YmGvM
J3XtPYNMk7mIAHhg2KyHaHjORVqugOzClz8PD8+bP7+0+3o5FzN+h0759gpNdSNG6yAbJhze94UK
uqeNpqIrz2LpW33Hw9j1R+RujCSKYMl+A30T9zM8XoIQDnG1APmRX35SNbMSM5vzLqwE2CtGQTk0
Vcs2OOLw0Yy2smvTh3T+5EmQvp8Slz+zl+o6WFyoqVdr5ME5teZeU9i6oclCSCmMeyntT4yAKYOi
HHVPiXqLjgn/T4cp+59AqrAvLXkwXqtHQ4h0pOyTqBPjlYp1eJAbXCkW7hUQTUbejm48gYhJ+1vb
nssQoCvyYtSL0BRRTTeUIQ6VhBTe++ytO0aJxJxaTNyr/BtL8h3qSrkbJO24fwXygS7ZP6C7yCQz
Hd5qHq9WiESLBR59Ba7yJSkpBozpru1q1PBpThvwPrC6MSY9hmgfZB3ramY8qjQ2x01qCg1lMTkd
dNaAnnRz40LNnERZaUJ6rOd5Y8Tj96c5YHVn4jkMCTMPcwCwgwHUYHZmNxbqtLYEwr0V9Npdm0IL
jxwLyKr3VqQxX9oRJY9KQGLfipgK4wdYvp/BrLuSUZUKkX63BqeHPYPB9/JJJ1P+nddY5F1HHcTb
Ev03xmTbQOhdFWCsElcoXiKUpY4UG7rOitfzdbVuN/XydZzIOPPbG7+9drGvNg61NUyEgcScMO8I
acFbenV5uv6dNJIaI2XuW41P9oamKj/up7V+1iyxdrh5b7viL+te/gD0xYR+C9X841QFRJs1Ec3x
U0xEXl+X0wD5njqZqVDhsPsI572IiTHp+gvxBnYgZiuOaXvcZYuGKtInNDRqaD7HIQGcFJIr75Ox
wriOIaJ6ou9KbtpA4tSv5ODXOYEqr+aET1/qyGl9SEuE/QzwpEdQSzfCRpSqy/Dmh2L1N+DqErv5
TPcL2q1HHSKhIicMvlLSRfXTczf0yJQmZxqS7pih897XCGmDzerzPfnb/s1afAqwAyNSVvZVj9sD
wQ4NUZSkzUh2XQsNYVFDDkqhyanGPEkDnCxw0IReWE3DNBmqeUgklMNq0D0/u70dLQP8uXYW1760
arzk1KW937TGlPE+lr2oP9B/CqpAaBCuoByKKUFcuUz5hhjUbLCiBwWvLXlR4r3B3s/KuK6BgTi3
Phb47NZf+8ojhtA7MEaYlWoLNa20h8uEIdj2eoBZsRsMwlyVdcrFxxpG34u0fvrhJrcQ+6bNRi4V
BvsTuD8sV/BgHzKI/9CprZ++ZnXoAqM51Xf1bo1BZQwb04AieC1ngPqFQXyJheA5JQyLCwak7vQx
/AdypkRNwCF4zXDN6TRu1yHR9W9ynCYYz233xpsYS+rb2ybP4HZzTLjILkMsBq9EHkopOd8HWYpA
WqVVJygJh1344JZDObPOAIfIs45RtnnCUKANvFdg2G/TG98FR7VxCYMqBrECyLUxS9Fp4TcOQ4Gu
A2yQNl0K5nkV8DvPrjqCTpaB3kqWZQxyAKDL8kUdEUA6Au3EWjaascm3R1hvi2qa6Pw+CYvxdv5a
CnN7mq19qc+89n9ZaNerjOJKDJw2xSLZt3AY0rh+VZOT+P+S12xdPhtVlOsWnvxZnNKQ7tnbdaVq
AWMcvfJnOVmLFtx20zeSj5NSWPuM5Rj5WNKfp6UtaeO8DNKhPKm83XDeYkHE8BFmjMNHAONF0Eys
OSQVVV/HKmYcarnpRn+zSyKbf3Nwgy16/u3rNztY2vtMDJUw77btMFCsnqbDYzs1p/mQGpbCS1Nt
SxBulGySfJdGJz8Y8CReJeSXNP0Vt4xYWAv48Iplr6FLsb1beOIpQHC37vE2+YO9QO7UCJuU1Frr
sbEwY2yaIhDJJKxP8zTNo+uEE7uCvydtCz+6t/YZeq4OTX7zZuLAnUcSIhWooJfB6oGNH6g72TBF
FrXjPYU1Ls2faRsMnHVz9LQwHoqDHMGhqYbENnmxPXTV5dqsuqw7DACbcyC9/Xs/5vFK2Ne+eJzI
5bA7UaQ0MWlNtV/7ELi6zV6hteA9rF9eU18qPh8z414NlQCSNNOY1/foHnPLphB08zGEnmlQoQva
TnnqSRbRv8RpEEiUfxSSf8xY5qsx0ixVUoV9Z3JaCY2NAZrTlpEUuqJC4qjUiTyaJIUjLXpcODhh
JZwbVooVUlePnkRSXQK2RvxMrmG7AKKCD846g+vbiYbagce4H9RucemdHtlE9CiFKnxfeE7OauyM
Zk8IIlyCdGhwQ2ydc1IyUodqnwGWTegig3+oOYwSLA06Or8lKm9hcaTyucDG5uTw6clbWCNHaBCr
+HlaSr0FxygiY9+niJmjq/gGFYxGbdnwbOpH7Nz7IRLLJejMehDU0K0QEiOBXMnJc/LEaBbxm958
6uiuVGA9pbKxfgnB53px/WUv8mc3lVRvnxoXwm1OYJgJXvpIVwL1DnTei0UvVRsc/8okV8vAPzDg
q6CJaPmXMTKKLj5EludlnTWVdoZV5xuBlfYD8SsQWTr0rgZ4s0KsKM8VaqQRxn9iFQo3KWvk+ED9
snVvvi9Zp1EE/gnbgNGPdOPIQUl1hg0kNnfYRs2v/a8PTnHScaAzCunJH0PxMRhZVUcmm23ON694
bJDBarSk0aSE+r8AtCFtk+rNSfNATDZYyQhjiExPd6lG4Ybko9evUhEH64fBxYPV1+lozV02wPt6
/v009Zr9ujjIIcSl2OMqXtrDC0zw5is7Gs815gGK7i0nj03niYySVM2GE0bl2fkXFtgbzpMQrHNv
I1sFU/3m27FXfLuz0eZGOM1jd2FtEzAlcs+H3yxEYM0uI9+fCmn3H7lI2bCOzfm/B0BIwy36hp8U
FOU53Zg14+16VIcez4CIa38KiqacW5Wsd6e5ePuPsjZfq1fTDgKZdVfKUa5LvEJfP10r0po7SCFe
74x8L/OU0esoxJp1PtePb05TIPcNjuyDzcN3UlBG4OOC9snIbnWKO/6Ldkd1N+LbNxRedO9ZZPHg
ipRCSBL2nLl++TJZSYJFIMNDnn1TjBtl1xnmf4GD2sfR3LfB9OOEue/0h4l4EAjA3vUckK9atDqe
QyUFU/r18x/FwZqURZyB8PDjT/8u7LLoLUwNwJle/2HCHBDfKP91sMJSATMs4xW/WHYEkbalIQLM
IE5dCR6kenpv4O/6y7REHOXCaBr0HU4W/qWw4yv9Nn5RMOFZthoRy4l8JJ5+Sx2AbpCZm8lzgrYz
SUsS1QJPOGCHRhzr+Eh9DA1ADqCukKvl2PeSxVGLD5CBqk8acMmQRX6zDlvyzixbD9v/JAj/LGkf
Pz8kgzgN3ceEvxRJj9N0jLex2TWepFUoYLWq/PBse7eClq9nWnj3F8yxXYyOzeHbxFUchCw28RIC
Yu7C9dsnFgOWsxA3wUUN5bqXxyfLWb/zwrcHjxIJrS8gL7+7JqgOVDreV6tWRKquVCnD+nAivDNY
qErAwYZWFsoOw6ye9kEfbNUG6yaVvj2nYkfF25CIhdbYkO9QkqmJWMbOakoeXOaeHdxLumkvL9eS
nutsHzWsnuB3m8fghpSxZsv8ITObuN7rRy9VgWhVREZ7HPeVdMmJPhJUOs0benWWegqrk2o7UURR
HHpfjuRqaaTsjgwgFBeSQmV3bu8eXlpaluMaiN/9TUuLrD+wzyeIbg8Lq3ahHUC2hwQQppY3qaVF
yiVcBslc1lmM1y2/0eSTNWHKhFXVzqsofJB8kG0sRbMIGE8ei6MjgJ8N27fcs0WKxAa88TZaspy/
d2T+8UM5ZPY+YirWgxNZY3aOuNj/KpJ+ELAB1xKr7AAUUH4El9kGEQtIHkFhT1GPkqZrOPb9fk77
5NZvt8LWp/7BkMEeAGXWQuYXmG3nZR7coBQ7P3Z+qJzWym8qxeIpQHW34l0eRRk88pg34LnnG78A
kSr/ihqjZg2HCd1ZLfyaJgrtQOdbrIpoprAN5pWHJAyVtjFWYeWMIPXEsHO9Gs99X0lG5ykymN/I
cSjzskKKHO4GqwC8x6sMktqrdf/8FR1cb9HQ+bFRSQYrvYiWj4/HPJ2NQwx4Z20RCIaC2w2xUxnD
aenS2xUtIVbttOhFsTFHktXJcpcebVJGFUWtkC76VmFpNtSoBpVWhy2v9j2SwJhzdnrBCpb153cz
vBlUX/YTvGWwZEzqtfyYlf5J5d9V3VG2Nt+/98ABcgWiGXOHukqsPTBI1V3OdJvSu/F8OAzuZqBQ
hmkowXqpI79WD3jy5EHuKfj7NOlBSR6HhmNQ5G5oBQ9YzfvQCwov0FOd1/OuetMIfZNG0TjoK7ay
ieH0njPfHfHQxmXuQnJWv989tUC3mFmggX2s7hodupcwRcgR8zPCyB8TfIpn22Vnm7AcHJfaqqa1
6ElH/jR2lbI74h2h0n3LhCl3npB7robiO6jUDv1wbP20W8g5VxI/cVs4FEbZo/sgN0YbTguiFCMf
t6GjLcw56U1XkksdbbHakYBevZitnAbc7Ho8Uhzq8CmV/IG6VsgdgK9D1r/UamK84YlMRoACi8i+
qMiCV1DFIAXqhlsMBsCVRfVmg4ef2nuI72sgl6enG8q5ZMGdo5Cw9qZ1JtgA2WhD1Wi5qowF3JN2
q6NxLrRvkol08FkLBoh+1li58/soQhVTRECYI4hlKqWSMVjBqh62frYhJjLd3pSwRl8MuNiiqdyC
/gW3S9WACLigzeWgJiKQ6vegzNwhufrE+VuM7SlxooG328O6oQZxvi83aQ2ep/HdrNaGLCx21q53
aCnnkr+pUhlRoF6QOthlZqM+Q4eXVYwbKtquUDTJ7I0xrIYVVLBlcB+oosJSSJwHOCrvRB4r2SLA
JsMMI3uDqDOAu7KUEfhpZwUrdHyy6sPYhksjmywBuEa9v1/BlcCaBpTrUgXjdd8AwIKY+er7ZCF+
Ubi/zkNm2e173MUL4qRCdAzrRsKxSlNQ44BgNylb2Zv8MzVxaVjfDIHSz23sQm2/jInS4E9H8axL
AC2QDy6r38YN2LLjt2/kw6sJpExWhjsPlNTCXgFKDlgGTNICumhJZ7UYLoQmBZUkoeYsN1NtpFav
QzuU7DGCWCcYnN3q89AohTaJD+Fv8aK8nBZVNe9vZsvERZpYUY3DRSBIJlDqJgxJawnPMTyRPl9A
jCV8BzxCld6XWr7RuhNPviIp2cUpqsaOLM96qAYcukoEJVVe9ili+6c4xlpD0kNDTXZMxwFO2z5L
7kVySqmszysyzzF7MosXReW4vGDr/IEdQvZunPwwbVzdA4UzxmlVoSH3DT05Aaj5f8jamkqN9Ik0
D43SREj65GzxfW3Msk2Bm4X56Ln9bPJP86/kRFkaXNC3ZBzmUzbt+QRtVsqi69msDHf8sBJ0Fz8n
vd1rI6F9z5Tg8Gyx6tNymwP3GmFWtDzroKoXP/LoHEZuCGyOL2k7pb4sCvpycul3wQuqyXlzcXQL
4twYijXmrhuxme2CTwPw5qJ6oSYu/aziRQiRhn/703vQumofM1eO5UdpvXdW8lgEhjowNdP9G6xC
jR/hYu5gz7dg9hXWs2RR00DQ1+K2buXwZn/spG3N8ch+DQYUzi65h3LKs6DIj7rmLUvDhyWSH9S+
txuGQ9cmgu8NmcVIVzI+aM1IodxDd4pNQlv5VjjjLoV4/e2rDDFwcv3zZLZ9GwEj0ojPL5Pjz143
UR/UgmJ7LrPVl/BdAr8F6ackkAe0Nj7POq1UwGPEfu2/TXE2mRmNh1RnGZ8dZ9b2HfSwzK5D7B/C
zhJDdpW21szTbpHkvhA45g4b1hSmNi7hWkR8hwxWOd98XpyMxvhBA7VB2gtVboUfi7oZf6mvWllm
3TDss90F4CohQtUfUBwqmyhH9/25ZbWvpAyyrCTSi1oilScnwLyEdBjYPLiQec1cUXdQt+f5SOUw
LG4zbRgiRI3xQHi7gt9tqFrLUz8SXyF7agMyoRYar9OeW0+ScfysSfcf+BOk60VgEwyhkSC1/0yX
+oDKe8CDrtwqqkD2WgzRcYGPKTeJbzlE49zI3wPSKptlr/rfGZZBYg37gC6kAgSLAeFnNj8rAh0r
Q50xUtWpWOD5KFQmck9hMSd7wgPt95aQJM7Fa3XvsSBj+JwqAmXsaaYv5Gn3Cziuvqky23gGQNjP
gguwXQFiN/oBRpVd+PmcnPgLpF697jDULDKGYL6LdpOiypgPfar/y3xGNt0irfXZVTJswY1Cj1XN
aNKT1T1MhYV/Sv7hwySjQTyR7Z8i7ESFNj/kwhhE+EVNhuRz6OfjpPeryczDibEScw2+Q4RSNOF1
FWhcsKEFG7dMH10/nQEtUd6gC/Z2irmWWOOd+cKXhDtMpmHYPvETT4lc8oxUSnJ45FovjzpjY75o
IhZXmkGzlmB1EGIx5hrdwapALQWfHTtVAamGlGIkH7K+a8iHaT1a1G3swDTFiLwRch1YP/0Hmhu7
8MSro4ShcOAhI4IAxYT+4Y2TeEhfacFmcH1hsQhHtPwsVi/LcUmoJd2PjYR1CebOEYm8t+WbxeRn
I0TA2lpq2qBuJsJyQ/F6IECdFHPFWBQSmgujohQen+X9Nh7Ahj21BKteC3KPJhpotdXPuwU/ceWq
73oX+99xS7Qw7OIrGCjV0GbhGXjy+PqNsjNfPbVn+bhCJ+cqO4ruarrvdFlcTCuw4aLIqnCOy11K
UuB+PM3I6baWLSVuqlp/nBuyNjK331zgYUDYOobSZuN2xHHDStwUhRzpIgJdEW+VCk36y6CjW9Ld
YlGJ+ZE7f6oHdhgmLa2gRL8/UNZdMu+giU+5D+ZtfuY8u7rfvn4dOmfIM0wMpGiiJgQ7CLGtJIvD
9I2Tef6SceXf2r0dPsDrUHckq7AGp/NDdLwxJeOkfNjx/cky2nAaaKnF4ZggHG1X13r50VstSTz2
oAMr1N3dZkIMl5R6HmHaDyY9s/QWAc4xlkD7DUXYRJVy6e/HY4D5BjjRMP6H7YF4b8D8BitFdlPd
mt7C3y8d3edAwzGYgbFRWZbpjxa27a+qmvLYf+wy8LdXxKZ+og5FIkmubkH35zg7jriibfcnGDLS
b7/eItck4NnVk8sD7o/f+AZi8qHgm0yEvuS5AqcU0stewEE9v71xyCKCFufnKB1yBNR1no5Ga+73
8Ey259PyutS0IZziK0hEJhaw0AhAiXaCF+gk6LOsc9zUYYnSPky25yL26LSfoa6TYS3IPA3lRZCd
+z3vMD+uIQ2qE25m3Cofwl6Snzzme9khVPmxmZOmatbP7EaJgQvgsC1dSmPGcKH1DvYSrE4IuLWi
Bvqqy5/r4scOtixmkbRCNQAKgbZCc/2eUpjWWzXSYYGNPCdYXy6QIH8eiX9q5OVptqY/6y/GsSie
JCMSSpB5EaBPL/7Y1GrdnTcnWYzzm4zS9dc1PwcwsxaVWXkfLf4X75sncwA8WlVf6kaC98B/pBLi
jMQqNmDJxWtZs4jsbzGOA+/EYEfjDbA9OZh2iQ0lXXYx0oue0C9rCd/808IUqG+0C4AGZ+izYWsv
rP+C7+FP6z/LKnRIhwPX+1hsRa8eGUGYbkrsttajun16R2lPFbcIIGMH4C+kJkraOBQ23LyFl99U
FBeoMhDcmRn/t4PhgdGhuXaFgbMHEpJjjbY+bEnz5hT7CF+pFkbjMU7NbviOVgFs7ZjMFX+YWywU
RixGmtGKmCjtzm2uJuzmXsCc9aJpVSC5w+kc0nKGHuI/WdEqnlDSKRNsqv5LKsCh32mhgJQV7stw
uZ6sHQHJU9Hmgc2fG2rh7ncdDmBqMLrLDDQkoJS60DmJAI9jyIsF94vwB3FyLeF3WSqo1cBYvPD0
58ubRTmR0B2RmzECKajfdXAZhRDTn8LjFfON4ZZFaQiGS1cLt1UdAsvPvvqvSTrs4HdWVZHd9eam
PGN3xHna8TvnygibBvB/DClRVNs+D3XQDdSxZHDsO8OoPtK5XaIxVD+I+UadevI19XKxs5AcAAcx
O74SMomZf/lBxF+eHl8PExKvL7hNnbVyV//CJ8NqNh/3dWWEpIMG/Y1fej8rM5zvR0DXJxVXSgN8
e2rtRU9FDOR0t7CVWSWowBHhWiWso0iy5sTdYWharMtWGKBe35K6dEb5oWcEQpDYjsSpbJwpAF5m
jwuP71Mmej+jMAQhPI5quf3VEOY99ACsQJPbib9m17gh5F8kWYRQ4vN5a+i9HGbXfwLbcwQxvbJ5
yBvEjgQfACtAQWL2Na/CtTr5g0pKBpjuaZOOS+McH7Dit72jrceZCt72bMPm79vvXRItdyJz+myP
mFgbDtlNzA9tO4LjU30FvV5vcKvySro8DZ7JuXUburTidDGkmjUa6AFg8WYhPFiGLAC5hZBIrke+
IMVxYHH2C6RBM6ejzCOq9VqKAfaoa/tDAImvVbOv8E6JfJJ2Blv5jip/xv8YbBSAtAkkEB74CZl2
+pdLrHwJvDsf6DbbEbaEFRbvimMKfqZHSrvGbsVvkLhY2W3x8tu9lSJ8FmNygJQrNIgI71BOi61m
+73C0FncPbNZCq7XaE/LwL0+NCpUAILOo9YHeNYrdzlJZflVZ4wdxvASbjNub9G3yitI5+Rl0Ve7
K5IZZmGqXlMknQjc/sHIznTz3PL/wTA2NgMivFl0JHFIk+5+UTOlKQ8tlBmrTUUbISyscXn33yNL
UwbYvr5uKIHv7nak81ECdN75t0hSXEnVNiZYzbRnPI2+mTU3sOlWHJeb4NFbFPTMULuaL4jYhvzv
xmdmHn2tktICxEh9vK9KV/vIwsLLyVPnwlqmNqlcNQiL7AVVWOdGrrDeh39H6jlDYQwN46WfIo4L
XJL3LpQDPoWT+yrT9i66z3efDHlkWF1jqmHhRT+uYikisMXsrOg5LHUx2FbgFAIGN2x3Uzvt4cQC
3ppsc7w19pGzayGRlqbYsGIY6Y5SLZlOOgJQv/JHPJIM7N2PiEGcdtWrdKj12Sx7ZHxdeH7SKkS/
0r0o7AqJNb3MmVQITbh1PSrpdD6uC8sQbW1XFo/2RJMAUu9F/WfF3/FZPGJITjsnfBdOyvOQNgx4
RSpa/nhCPx9Y58ECSsUIeLQjy4qrEGfTO6jKFNRT9VRqzGEJ5aB9++FV+JQ1SDsDXk4dTbTSbRKj
BJ9gk7pnMZfrFiLtwRnxbxKCRPzYw/zcbXM8rQ3kVAbPjp/nHXz23btwgpF+EPOEd6FT/UefhKcD
W5sJF4GED5i9NerPFO/2L/pzgJ5vH38olBftO5nBk6Voxq5yGNGlH+G2M2REoNmefmStrGtqi0jA
Pd3iJ+Y//yBqhjFyUpTz7u6kiCJKcqYM6/wQyh7nY3g8na+aPZm38Ulsi74HBihH1CRYB3NbkTKZ
AZLYMWshTeiQfXHcc5GYwnbj5gkbZmCn020LKjwBq4Ag5c7Px1+tbDs9OwGwO8al4QMUL5A13ffA
WjwfWfLYH6GgOAmgu4HN7SSowQijJ2mAx1CvZPM0bNwM/Spt4v/2XRV/Iqugep18+EbOmahb/O+N
1jn9E/92hSi28F8RtEM9urZ2ywksybR6qBKduug8tmevabcua7h8Uu4L0zrd56g2mC+PLOx5/s0X
vvQlWOVsPSQYPDx6kpwXbuvv88+hxEUoeHFWurdHafpdBvAzN+w6wb6NmLmLsJJLhNEwXSyj6SYX
G5bNCc6UPQnnNeUgLWlkTsPzyQT7aUXF+PAGHYDR/6EPfgzjERi6OTgtL2BKhamuc1J4S64sHLxB
fTibXV5S7rhhPEvJIikvySdqWGxMnuxmhawXifSB26Mt2I62bxuOZ03jh1/1k1ZnepxZh5JW6+1Y
1a4cObCddGLmMqYadAWikuOhPK/nyC3yL030fZqJR1YsNRoqmzNBjgrISQhxVCNl7WaO8KpHJTT7
BCUsEWRpwTY7U0vjHJH0o1WgfhLw9vpJA27HAEQbU9yMgBIsT/IeXLfYEf57JpHGfCVfD8HIgmiW
bXw9/IisciFc1gh9RNtXItkjPodZmxQ7Cq44umrnym3gJAdVCT/jBVwhmerv87lWcr+cIvBKuHH3
+uQDJJsMkLh+JnPkX8t/43suqaopzhBqH+ghR6x9GA6dP0EQ9FsMAd8uoJu+xzOoWK00h6DDuWr0
y0oaDe4/VyHXIU3vgkjPYYn4k9JGTYaIzrgl8FmyQAgwi8YetiCyoTUoJ0nUDwZZ4YtcgpEyavRQ
Xx6WUTdusA0LrV9J006b7Fl5NgzmvR+XyUywIdtgZqsw4TXlO5DTsttknZD6ao5HoCcB6kUBKwEN
ZWKd9TPpulBq0xFsxY6eJnwKkUzEgGhltqkP/yihtgovJGuXiyf2sMBkXXrgXMsoUAYQuceqUQwW
9lbTAvPTF3g+Tq67whDSWNy9YLPRntT+/zGfOXJND8MtcXpRT3QQA4lutVgLZ7V90+y3JEUeeIUM
c0t46stvhrGtaf81hmcb9K1AjOwXZyRCQXQQ0Bu2nfcBvLK+JGgIcW88Lw7MBRjYM9k0+6eZfK91
lkpHbXBlwnfK0Ug0y8YB6DXhHjSwzQs14P4F6BUsmw+e54SRrZPWO2OITY5HrddJOKMydLOWpzdJ
zWs2J29xTcyooweFKXBOt3zxBilcxuKUb0dYp4FzFkRlIKMOg6fwalivfZCiQU6d3UPHAFITjxPX
T198mcvkMt/EHVApIsP+1QoTaYZr1T2ks9M4h+NMniHZIXo+mOmwUAeL9GJcWHx5DCw9zKJHRD7G
U1WgY884KdV0In62jr/TEE4ybggUAd/N9hjsZLp+T5YjTU0pXlxWLQuk4P7P4Ui+Xr5Kwl1DDT2L
MHFjhYPDGK2shCT1Bz0sTu0dp3oPYgfKWr3X+wGiPa9wzHPq6AjG4vsOWOjMFfm4KbKw9g8tN7qA
P5YMyQ+23omayuoy5Yomw4M3PrAyzT9fGBi1jdmPaeoEWMn4y3TIuJNccLoc0+3QgXmFXJrdIS3Q
se4uI6lmgqCOoTvsZqpROazmjTvWFKXuV1xYO0KxU2D96j7r2eldLjC/6A+bMn1VdYS1qDRJrd+r
k/WUUmsWajOIsG5UYizkeCyI4tdnNgR8MEk0Amj7Ad9N6pLzEqtY3gZTlnWY+uppKyZ5IQN6dQtK
jFbdeFJPupYcRaFUyE2ThNzmH1Qw8D4mKgf20zKkYnTS35j0+XCTiMQz+iCXeZbHXjTVHJQcUYMO
HYLsNXTWpp/bNsc/RbFDKfVaBSG/xzrLzNqPBhmPtDHg1In0OEN7pq7kxQxCDshhTdgq7v7arWP9
HsiVlSBwkLVfbSz1OSQgPlrpIhD2mxurumNirUV32wgg9kfDqzVQIkM32VnNSo/RhLC8CU1U1JFD
2Z5nR/20ihXLfInB+8cbuIxthvOcZn7jQjhYn11V1MS54rnnFadX2A2m16gfvh0wGMuS2dqm0iN5
DSEFvKSyoJZnhHdojh30njZ7WDt4wKZknnLq7pT1Vlupp9GCE8gHbl01s/N7PelHfD+BX30kqgC8
ftjZ1xW8nr7zTG0DHET9dIP6Olv305yLmwArMa15CawzmvHuu2iEajRVXqACdh2qimXx87sDavwT
qLiaAb6yl+4NDl+9aOH76LzpENmuOxod0U39VT34Bs96Zm3RllqpwYAYUDN4HRZnWlbTyoSpJwcp
9q2M1nH4FNF/SvbnXN8qs+FbUrdI7UFSTTJRlZIwOZEGBhCjL7/X0agQIoqx/x42LRPg67IuNEJm
2BHQTprpfe5RUxP1jhpYNSB6E7pkTWJcFP36R2kIfLO2XLjCetY3J+3ZhtZkHxGMGfP27gYFjrWd
abnT/GBNwyHY+ixo3eHsC7tyPQ9y/0B7Qk/nsMNWThSZe5CB+cg3bJnMQIlCWAX0EVpDHGDoX+vJ
DcRHTsl/5XUjUVmiPu5ZHDG52uOZPtbFc3FB1A2dSu6jz8iGye6EBy7A5B3pEvxos+qsrOdtAlox
GipVto7GfiVfHeoNrLFGYTN2B9Wn/sSI0JM3RLZw6+ruXClE7c76+psJelW8KOfaeb8gWHiAzRpf
yYGm727pLP8BPCYo8rgTZXYgkRHexFvW+4uV0Lzn5vCxWIafyNzSsJSEzsvXee/6PskIA4wgptON
QCnW48CiT+QZ9NK2bntYvl17qlOiIjrgWj1MaCLQo+K6HmVUP0XtUc/vB6I6nJwryJVqYnVjN/rM
6/yk6NQoQwcTus9AT6gV+DoRI2j0HpJx2j8biJyGBMlyN4aGwhPQnhgQfOtPaeAf8UEBocOaDMUb
aBEQgKRPEMCJM5pxK4r0cDIogni/to5dh0uFEY/iJtukUhq1V41DrzUPzSYYQm8kOjlS7qmlVQkI
cOzFexBBzQLIpvFetm4IpwwFDLyqdEvsIJTSMG59YAgqqWO9yI67b2rbHj390okNPDNFa3AqgzqJ
2MaIj25mqhPlrvmJSTwjkRDvsKInuq9IEavfRtvFP5H2KFaLuR0JA2aqb/HwbTrX2zEe8rT6Ti0i
07OE2qyDyQEk/VziFoTc5e5isvCvzb955zKKqn/9GjRQOuZEB5ksLOPV+ytLIS3H0mwteAt+eCNQ
jZ+ahML2uKHcWKhCn5dTrmq7Tr2xMj7UOE39Dn37BubfDtf4lVFJU56nqp5E0+MMy1xH0ij/Amq3
mzGme93L1PUWQvdGVqed8NYY6NR04lRLQtAqeDUFziCRhEiqu5H2H0MOMCFGhkWFyJVCn0YOHuta
EYa4C/JbWnK7HpktvCebS1ttDCS2HNPtfxXhMFV0b5fl+KZCNxnWGZvzQ91HJC23yV7WTkoNB96G
XOu3UCjMXgPCXo6Gz7hPBPAm1QQ02N4wAOWraMseE1zsIlopIppOU3wsfm5mPeJ/crd2ZFlJArcc
ofi6zot6APMwoR15728TlFBL7qahOEmwWUGrqxvai+LVD5vUubmWp+IqwANWMD+EssxK7drbaayj
xxDbF0Ehfz1saIQyVZUsz+uAQw6eKBKpguG5ZxIXwLzJ671MUCekFEUIldh8wEj6PWU+pju3cFPY
cGY00pclzSxj5aIBC4CDY8aQJDBiAUnxlEElif53OrKpiDXr53QCjao3ok/BkU84yR7YaOLWXdbC
SC+oH2EHlK3sTY6Y+CscTNsu5Uscj+iR3uIKrSOiezMmpmJqDq3Ssytotj3O7pBS9NlQCZXyKEYR
RjR88z8gA7iK3IJo360tniTyTFyEgufS6I41bPNUDZXqUsyp8YiOUnagsgQ3P48KwdZuNi5YuOFM
9LBV7QpWrM7VFB0qdWZxZ/yW0dGp/w+GZ5/GJbvGXqecXRdfYme93SFRwTShd26eH0lwn9W/e15g
mreZgFGClIwdp+YJyhpiMaAGuBCW90Q8zbGv/WX+HW6C97cZdQOG/boNbtvnEk8sQxDpoao6CufY
zHLO5T5dWZMft+Dw7u2IxQvSBd4ZjhYZ1JQ9zMIB4bbABr+DYN6cTGMw4e8HUvrR/8+sr1n2nb4t
Dpk86wVI1r+V8rVCVOvZSX3CW92hkuaeRl5fWTJvBTc9QR5V+Y3bD4QVSyuShc3X8/sB6lfF9J0U
hQJTB9OFhreLKl65VEqXTK9DivzyjJLSV3zXjDecKokynnxeNaD7k+VJGD7APwcT6stTtcSiBd9c
MP48+4k1qlE/aMqsBgIlZtejfpjx/fXREGcNqYVPOD+u4JlGDazIj1BrVXdNvShBerFCX4H/guSb
RjChjsGfCJ7UoMjYNy11ciYHv1xcyB5qYk6c0XfhVDFmGxU9Pi830oRYxa1h0Kclf+j3WxpNsIEu
IoI8VGjn++/dMJluhz71AKzNqkoIjXEonc02vZSU3YfOdWoAVe1YFY/pE1bWpvr8bejIj/YJHHSP
a52iJX8Y1L3eb8WOrJbahrjtfSTWe5IZUZwsEbGa9/HMu3bpvlDsR7jEatFVk3RKCtFKq7VcJ3Ik
/wcugN0KnzwFcdPH+4cBmZTPGcALxTcfYnRQ8ShB+erTpcAryV+T7DfeE6n46w44fVtFDJ0GDf9L
OvLIPEjCE2R2n3pRek5eO4GOWpl4THaYmRcnSC1fvBgTYSLWOz3k/BLSzVYpPjG4D61RpER4rVTv
uuUbwz2e/PVvmvvNjQ43oE4F5SqzavGQuv/kkZMkbmMzieT4nTih+SaGcroc3xblu2CAjAcA39F0
ROhErM4Dtx+sj8phYbxFD8ol2E+sbyhyrsartPELWA/+/P9MIR1qjwOBsFTp+zEXTWIrx0UY/mDZ
gH+9IO5fOnES5b5Bdv+fekruifXlz+kHZjiObeUO+ykZVQ4YWiviKxkKWYgtV8M6w0Q1Mwy4484w
AFzYg0mR03xi7u+VUC9mZmmQvuXBKohf39xeOEXtvjvi0NxTr25zgonrWRuo3rbqUxL8jyVB5N0x
MOiqyF7wZ/hT33Ri6ko2sMSToAAFql/BhU6EA+1l6g+SMT1OhEHyl2v11PtvksgpuKq3NhMJVX6X
+zZ5XK0VfYG4ZOglihCbjneexdQgtMD5UBtWOrl6sAxo5sHLR1XeJ3IkcXjgdABcFeesvhRyy0RI
56vOIbIYvBm1Kf4xqcTJsxPR8sVxDQfSurYTaR8gTSRZrfRY772XwFxHMJQOVqaihwJ2o0RV+vBY
LNAnKVJsJ/nrPt/sEPHRLm+dYkrHi9Y0p3k8YPKyDQgXh8Aa+nERvrYoxikgkVkKhxrapjxgEAf3
+u/HCx4pjc/aI8FeS4Ro/t4EE84HIhZ9J2pCTXEqViIFRPSxdMWVWP7PVPTNz9H5IB5lAyqtTzLl
APxiTStmJbaXBeu2uMO1jmDdnAOll8vRWhLGkSZqsCj+xLVG3cO9kiQDKKQNWXMqGXzpYf3kh3LP
ASHkk95bvIJoklHL1VOND3zEPgjWSwERW5oCm/wOLmi1PijhzC8GAsU6OfwBFtg87EVVopCXEHYB
RdPDLALw1U7XTxQ455tNvxOEclKMKP3ElRP7hXFWGPUxU3ImrXZE0MiP+5r9/td6gOabeRCG80J1
OHrLOF97ULUV4H05063pDeRgl6Yon3pT6SU7ygwJKbJ9z9CFmrWHnUH2844rmO2tu/0PqoimLH7a
teiRrg7IZyZX6NecdU1DARA18Z0RjaBwlEPeVPP8AH/HIFzgHbOai0Gn/wRpl1rLO1WybODZegfX
cCZMDiYI9YIUhVtd2ejr/jA48uMpNFbi/3aHHRfZGANrS94EATe1d70GlmNjx0wTkiPSnFrde5uW
z6BaoGxR6OKX7qLPFFjApBzFs71JOOkoQhM87utPJWwRAArAijjmwG3CFssd9BKD5Q9q0fwjG/Z9
qmjSu4VemEcdk3NDKyhyg7yMVfj252m+vLTaWD5S7zMXgOlf6Tsr5HJEZz8KqkrZxSpvcntTX2jJ
+g/8sto6p0c60ePVSoUoKMxpZ/Cpk8/LmaeoVFgYCAz2mK7qOEk+PuWcZFDoIOWaC6e4Jr/8XlIH
YWzfbQzxgNub4MJWVbkg8Q5M4IgeGKD7Ag3XFWqmAPcVjqanhgcqgWz+abawkuPViJLXcoNboFRX
6MGbMhb/YBGw0VgvinUsQNUlO0xnpf7FO/N3WbLw83lNWNM1gh8bjY7fyqkLfNCD4d5fg0FP0JjF
Sr8L1edy78I51At7M/HC/zQRYj+yUfZrpVV2ygMmwfsERbNKhVTofBf1MyS381fQwLYzA/7z7WuD
d29P8Ar5rN/Q6gcHNu7q4f3PCDoGxJdl+ZUMfk1RG0DKAqq0zzjhOzQ15QN6EjAOHkFlvjyEwCLO
wbwUVVRtE78URcyMhygu/kM5jNupquO4SqHNoJS2FNJCdOHwKSWYwxQ25RJ/aqdXBPyRP4LpLhnq
s2AJKrcCVP6ERspJsob9N7Fvi++lz+xdZADfuIXKgMrX+SIzebHnoqkEz4YaU2qPWzmXMyrkXv7S
9TVZDdAIah5UnjbU+PJBx0oiiA/qsufsm5PwoX5pX7RIPYQgyluKi0vh68uIfDUSiYjpaemP0p+n
Cg/r276hFmR2oUCghX6bcMd5xnhJ89Z3K/VB9H0x6QeJaD50fxWMRrONjkIbHKyJJDoYhLaK1JcE
bETnENGhnG0fNCVxivQVbVIUFqO1Kv7sF1XK5iS0TJakeoKGhJbfIeCjpr13vXvcY0yx+VhJTQlK
zELj7M3XCSz8S01XzawLD7p2o6cKeq2Fl3B1mozJPAOMxBBjB11BpxTGVq3fLxP7U/+dfeUkq0qP
WUhVvOsJOS0pz87NWhTdXang0pTbSgDejO1aAQOtQxzKrVOfgSLjT7sRyg5FKE9fj2tGjNVPf6ne
l4s+AEV44gOmcLaGQFVVDBbqu9S+sAymYM5nbumGfck/v48ce/hNqKoF6Aa6oK6sZD+a4eRpW9wK
WziIJmW3zKL+noJvS2l9nPgXDD7y9A5mkX+pHidY08iz3+tss/e9W4XcIHsJkWXNVTNjLzBy12qC
sQwXbRqaym6eGUVpZGkDM8FzGLYFocsYCRQZJ04JYKE6Y5Bg3HXaCidmbwKmRpNsSn9+yC7CK2k/
0RorsdY4T1mpHCBK9EEYb8tsrDfi7u1FUGREKGOwljdJNzWTK+RUYcuq1QEtv4Og5F1GrTYTvkQU
KH3GaWdBIgUfyB3EkG5HSZLk+bwenmWe6Dc6qs7BpBzLzm/e2zanT929dADqZ3y1kUAgHINOcOPY
/Df3ANqVoBgygatDr5lCj2p15M//C8PVoOGWJtFuNTM8VICyaj+KpqZsQVE6nalFLlb/3DIMkmDE
t9hkRfgfls42hiS83Se/EF8oiFQLWuGqRObHQkL6c/Rdogm5Ljvd2pjlqkoPva19TRmL6rqXqa8K
AK9RxrmF5UMjOPbWWSv7AGozfWQpJhK4U3Wehy89JIsPt2p4C1lgqp3aCXjQ2xT4xX1UeUUHEw79
6bEPY04XcfCnvaSbdmNZJCrpnsn8/X0GZn3IzXord8j0MdAHGLtHZPambEVAKj9cqNfkVdzlqKWO
+UxEoD6A3EtN7bLsj/kOe+Maaa054uIvWZDOYQLY0MaqVcP9XbXVpQzSdS5EAWxwg7R6LdMkH4Xs
jbDbyp+lXT7UsnOBvLWbGb3DLlzJbsVsv9W04inVTmDHuB9sR2pLIMrxcirbSBXaDNtLXqMDrvwY
dQPo+3pxIeH5JnfGI5CA/QnM9SxzEFA04Hkr7mv9X3ltuAEwpdt3V0arJjRCDg8IfSdHQ84C0Guz
4k5QjGObM1LLEVfVAylPQvXezo68G+/fllRVaBNhkmT5S0+hlKRRhWAbr+w7mju2DN4cvO+9IYRM
bltnRWyHUCvMLedraZOu/IrhhOjcUTHb6KSp76cnAy/4UpAiyDKgtEENr9PDXt8WQm8J7DxH+/8r
Jkb2kzeVk1fkLecHdLlanaRZKxVOkd4OaEWi/InLeHRLXToYoWMxcSLAgiWB5XHqfn6jVAoQNDLH
4SfHnrT4Oa9KvDeq+i+PFDBdrhfO4XJqmDidMMUY4LYMia87Rz2zmIhhADOHn2epFcGystRYYfr6
W1a5AbUrWQg1+p+dn3/0UAN5C8Y5Je4Qkxp5F57Ujhc0VoZUmHtA99cpKtcRwj5g7AwxhrrzxOn/
YxliJL018fSinrRPHxn9IDHtQMC/CqvjZOofp+akT8Xye9FD5zeE634Xui3DBUcRCFIbffHj0Kqf
4sipmfqE/8Xm9WfZ4Qwm7fBLRKSZqABBJM66JM/vuvNiFZ79vees7jrxr1mMTK8pTohdzOSTPDIL
9Ei8YPoeZZfiTc29TYsCM1+ROKMUcL5EIpAqDNyHTuBqtFBJG2nBVCQnA7ZXjpH+yKIAzBBUsjkN
dd59D/FQwxRjTh5far1HFpBQ5F4t4N/jG2F7Qvq3mLOlkR9d3sOeAHQodmKnC9Wfj4GOWsZUz82X
zaOqh8zM07+oMJLgNyGG30RQsddLn2BwdLnFGzV4oELe6swOJCvgPe2fD7RPFN7xcSlAdX+r4/wQ
W3J2iXwcJHfTP5cmDlFxkTEHcVm8Ey7+j1aOn4pXIRN2Tx2ZGNE21Ae4iDeZz1nPfEDtc9XAtpLW
fIfowdqC2/OAtFIPLHIw8fmRHt/9HaodLCVwwy17sdXAECGNQWuQBEfk3f+6dpzBW4qYh8CAdfbx
5U6vdlCk92Nj1HvQS0Yq3+1tfycKvYdFLHHrXJjA5QmjWC1sl9eebQdCuPkV/R1zNNeNvCnzF3sV
Tz5ERj1IjqW4d2gPmGOwrpCnIY8BPpmJiCsDmDlWedeGQv3ZnUo+5gUCnIXeUhr7ot769KTldNVn
fz8GBtDdeEWlSf9nUbF/8UUS1Nlhq2trNNpc6PFau88F8rYovonQYWLSP1osBisZphqtLhZij6ko
i9taiA+ypqJW6NnSevH4AFhBnMctEkJh1gWGlvUzzcAHpAI2TAxQ6hcVJZWUZM5RBymWlRpjLdGo
XeuXx/8J9oHFsSCv5zqGtdEXOe555HY+WkJkflPzHVdZIm3MKmrnHbnIw+QSbY+/Jf6oVuETdYWV
GmbGiitDf4hwUSlfRqlm3Z3afOeIilCLiKgMmO2gXvA9FjEaL8reud4JddgLZ+lRAUeKSQQqH8Bl
ZTYIE9z5X3txWMD+kLgxdy6ydeuD6aDnOLZwj8bK7LoM0Tw0VoDVQwTRRqt66+a+vRQ/gtoDVRmM
jydYEVizlBQEqzWIjt6znnU2lRf0H5kPqgTiGv6MCAYc4CJapdaK7AwuBv7RzsErALxOKeDJL8VJ
eHywsJrXIHHrnqzgTcTxW3snFKmY4mJURl1Pp7iLvSzbvbRIR2HiZWlEid0pLJ4TKo5VCs1ZOrVI
NAC3ZZA760Tg0JBVYIfiSv5qB6veXb+K4i1OW/alBvylsZ8sZPNntbft8a+L2cVIe59cuFxEy0NN
/H2/V9yCoQfXFW9LwPlned6x/Nr7jUQUGXIghh/bejWxBFfRMquX5rpBX0P7sW7WcBCmNCU4kTA9
P/5KenrC2eZs2hF5W0/BeWwISnABA3+Je5hE4jfa/bN2XuAmB4YltWcC1Jg8BkQo5RUrbZc3f+c9
36f4wDUdlsfjBg4pt34/GHRnu2S2ECaUn88U0Kn7XgMlDobvfa6EdO/Mlk6PC6ePfj76rE09s8aX
LtWYBqZI2nqYak3bPHK4lUtAQkuFzm5WFFW8htlbW0ROFfZqBJq+VD9u/qlnTrmG/imV0Ajk3g/W
+K64ZXTDvxJ0ZsvHpZIypxkHUisFQ40R9GQCws6Cg89R9vbj77D3tqFI3MnH5UcCSndGlPshDcbd
RvgeTRbtcT4VSqUwIHrMFFlu7Bvus1KnF3gWsxCjQrqN/BfX+hdTb1rEHNFGWCbtJInq30WMwivv
mpRgz9o9Y7vxeu9o8QPwqZMeDJx1cjC7QlaYxR1dqgCV91UUvRMp0k42zI0FWa3Cr0O6WVUWgKg1
9Y+1G1YMkeB3QeuUbc8c2uRPM+tfvKWrt7GHO3URy5/ZuyeccVWE6Qt6iV1PEpN/WHZxIkBYt+LE
MmGLeIYBVfH53pkv0lvXouTJtIqUvaynP0Fluig+uVq5aocPSi16/KGAgP6IpLTuWYGu6rOIJo9m
paFZ8H/feZYB7hxdIRJxDXJcr+7jPxmbcaS6TyT6FOH++DcpRZ4ZLQ0R6tnvfNFTesrc6hmahl3o
/SPJKZg/e/C2XpzvNYNrY8732+gg7ERNUx/gfO8uQQtHkm5RX72Sf2KXYl7F0gfYo7HH5yTjzbGF
1Bes7YL7KiSkEO76V+lzMlp0jPFx+XkZjSMzgPIbM9tMn5RxfLijSrj90D6h01NWBik6PI66eEfn
tG7DWVKR4dU3e2hxkvjH741J0fUh0vyIqMrICNA1ieR0L8Zf6lnAmE27vcwGy4xH1mfni3UG3CTc
es9ZpEXrlD85ajyK2R+OG2b8v2Ei8cZBU8XRuNctszXAlIfaQbyYry03CnetDT3ajtgWV+C8qHhd
raGoF26Y1qX/3ygauT+C9/HDGMZZA98gwOsQ9XuDchiEk4OFn22aOhMiW5qwqrVSSep5qYCPXWQJ
0nkQ8G9e/svLTx0z7+Df8XTUl/+HoaA1+OYv6Cf81N8W3lYjZo7l4cSZv20KePYMeRIOGvXuKuwL
IkAfo1kU2+JFq3omNVX2QXlO+yfsCW4QIOyDS5dHph/kgv9nq6CHJ8YkXjm+rDV2RJE2vRWNfKZD
f/A1G6zX8DEUb2U8WhZXLUc5zvXBZNmrUSbeLoqg4JrDwFdOPypA398bnqUouYTFZssOD1GWZGl9
bJSrVqCPdgPuk9zmmdcrDymJcv7lf8nnJvNu1a/f05EZCdxy7YdUCe/73NhnUsc7BSHOZ7wALF9C
HEAIEVYrI78YxBfCQuE4ihqVijDTMw1Kq6DWINSNA17XCVVUcPXVYO5Hl4azvJtvIaFtJTzEYW7d
fGAkdkfTAfSYRJXHBhoVM68xpO7GUwJnPFN46xXx8Knc/K0/0pBDp+gNa+yLWK1P80xda5seu3Os
eF4Vws+6gp8bhX57y3WfEHgaewvcObZ3pmVK8QuHWCKMGASlP+tLp18ut5xmxjGRTli8xmfZh3hv
buVkGrfcfsC/GGCh97RDt3C80ZqpD754PaYZcuShCu6wMwNVCIVbZpzBAtWtcRta8lKNelfWvFCx
djfkK2fVJi7Qqrn+2o7D5oWu1Qxyotbt60m8OU7qgv8efTwQe+ci57ds9iHBpk1V3LnzPMz4UKiM
EdCgw4OlckL5VN9ueO9gaBFs95ISnpA6+xiEFqvvY4fmZxF6MpTVwDpUXgPTYxIfL4l5TNQqhjJD
knBNBgDpqB2yHXTPxdRUvaVqm4vs1yGzmVoogQ8gVmqmQmyXW+aOUwwjFOKVUQRuaoBH8lzx2jel
bNCcVA4WOla7hJPKTJ6eexDzm+HpzT7tAJQeGlfF7LXo9C11yBe8jUJNiy+EVznsibpPpc+n2CB3
Qxp64TOMFmBBTYaChy0hyK+O9bN51RW4ihvSfmJF64P0yaCXWfp6RiL5Hd4UyP/kCqtzYWbJrS7X
MtHHruBWLXCXCe0L3iinA0CUmRhVIbLbAJc6MR/E4EhE8TNHtRTYmV5CNQB0jsJAyGktm0J9gyGv
KoGhZBWOHi7Fs4wi+ZDmWK7nXCoLX+jyg7jxL1tEaqxTK39GviIHdt8Xpl4hQFVJefw2nuAvg3Kb
x4wBheAaRViAdJ+3NaKreHSOV12gBIaEktsue712Ci++/uNLXiOVED5zPIRP7oGvFOvUsavq0GwD
o/cpX2JHvE68HyiaE9RjJL96kSmvHf+GfSieMa5FKeXEOVAEH9DYKknfN5UK/yyPvqzqXt2JiX2X
ZhoW5SF2HMz567IDf7LRelTyCSUk1ivgUUxw2TADAa5cJGK9bwLusQsUxXr/BWlI92mjYdPvBSS9
l03Z/5s/+t/CdBXGt0KPHvlyY7nUle/N1S1try59BcMetaXhZi22q5p3wx7qfX76QUBTB1tKJHBa
Ha+mhb9mp6+4KoOqDfNlehTnoBPr3W4TvpEPt8E/xrl6XD7/d7WS9M/+z5fQtr4DbfSDA+MLStmK
wN7Yd8cE53FiD0LxmVF2+eczRqRluvnl3Zmq0Vs8hL+iQajEDIDvYz+JAy/nBx9z1ZhguntXbM9h
mr3n8xSz4KsrBq2uM4fCZJ42FqRD3X1Y9MMsdynkJpmJmyeg8IDuEoG8J3PQFqry0g+vJqvzRewU
ZLrwxgcaa+vIX6fYZrr5mpqLSHoTLlW1N9pSLvLqUU100tlxDlA89O32PKSk1UIxMQw+D+t8XXPO
bHLtIZTlLUnYDTCEC5wJ47JS9vitwfaLInulOaSu691hF0cOI4VTvv9/RoO1RmjDKTQuij6h+CGi
OLWxwZw9JSyCiTQRiXCXKyz3pPZYkaO82xdqx22pkuEVNEshCmMdz6kgAAk1H2jT3YK4BJZI/vJ3
uXg9lZpnfK/wnDUwjyU4SkDehyr4dUHwLIz25a1PmWPpD2ogWPqY4HOIyNxFsJEQhgx/HJa5mfGB
mdxGCCqeLDxYjhvTfiNTel6mqLuT1SsUNGQ64cJn1X5UMuT62US2XoF3l8KSk250T8U3oHGOLgsN
zhEMMqOqalicVPD+kkQX9pdR+2fODxTgiF2ueKHoQW5Yq9HoH0xBpSCdzsD5tCdmaq45PHy6Nqat
eYvLaRX/qPKJ/PzH/yI/0cHUYCliMwwykhnwAVZ2KPO1xTAKwEr7k83j+YKjFZB42XtM+sw3b+YD
OXuK4pjB2rb1+V2yAUEH6GeBXecboT0Ke6xV6dj79tQ7F/ibASLHFPiINP/uXdaP6E258lN7nxaF
35DUgPGtr5SVdH+vhiYOe+RDFLYwsIjVkZMTQ4Rwafm4gRKte+vEw4XFafbMUlylAi2PJuf9rFDy
IRcQ8e3b4jYY8fdbe+UQyUw84bnWfb1wQOxJpUXjWBzNU5uju62zLsBPCm4/RVcxCdrw1e63PAhk
b6KcpqN9L4qFNpdilr9sR7CzsPZxqr3njRbmRH8i2HKI8oEFJi4hZ8HYbYGwaeEnqKUacL/KB0Ip
2Vwc5Omx2Jx7NeP2DuihZKPiNYPG1jQa16MLmc2iY48vdz9i+uE7b6sTctgUGPWH3GDWrAgyss4W
FrdLrvIMGZFVDmM1oga2w9eQl5Q3M+sTJ2PlDq+OexR6+5TTf0VqussoJyCVvpZD+UfTPP9vlWJQ
m4c85ninkUGdmEBt0bt3EzXDcrB/DYxY402eKB0k1igY1bKRKXnRMIrgT7vhyRIhcDnW1Un7CmEk
m0D7+IAxCSfMYDpby48kyDttjU1scyE8Dy1W28Uv3L7LKs+VOgZqNZDk5UpXug5UHMiy5uHbIxO2
rZ7HlrzrWNumxdnCVSIFjTDGQhlVCQUcCGaOxnDnwyrhMbYrCgsy21VzkWC8TUTz6sN/ONtCrOLW
a67tvYYQ7mKjc3rky6DXvTDzqlo/aG67F0gKJNVcZW6Uidpgz9K18MyPDS6z+y9SPmBH1Fc86kiF
uQavQoMuAd7cswfeyKy8WdDnhLImnDzf4alp6/yUa05rvAxLQiR29dimW4odm9xv6RFPhPQiLk4w
99o1qaNpWl1v7A6M30YQxqU59k2SoMzBS+zKrFAIV8LCtDNnAZBE0fG/x93qtw2IFLAHx1fBQmCC
CF/D08BOXdhgLD0o1vZupR4513qmgKUIHR+yGARAjDBMa9SGRiCcglq8L8EWWEbx2Ro5hkEiffZF
gzgp2ijw1g7pIJukg8ZQjBYOjU3VQwwJIPU2gbEpRyjBuPDJZcsVKxYc4K7uup8A3CvGC6hUwItV
loyjcwxnUYky1ORuBWZvtriZ9OVaF2GJuY92YOXfdDMPnK1RPomHikpz9W7C+VNEuoqZJVXKj9qG
L+Sbz9swPp82eQakPUByA345Vw7Xtb4w1R+HS0bcYpAwVut67P/q9UwyWEo1gHGWky076Sk5XAto
riJ3cQziGMFltK7961/TBgIMhWzHa8B9GBW35m5lwSFT357QT9Mkm6hohSgui+EawU1Ce0LlKar/
JDJGvdy1rsefy0BImOS3G16vxZCIsYJv44zmpciPIzMhdYFdu8W+O79cTv7Jp6bdpyyU5OzB8l30
Tgkel/kMXOSqV1T+C2PcxCG87eW0JLd44d5oyfolPzH8DBHgZyGVl/X0xAMfqSWdVHFdcYFI7yZl
havSENwWADAGmFtyimitN5gFu48LOCX199nOU3noxSxA0DiCssaAKLgoDUsENFpRwfA2rgKzuKPl
VczXbk/FP1SHuZVEduf1aGUIbJz9gMwM+DGQgxnM5KPqfqzhOFzLaBElOe64sb9noyum0X5mexNr
6vLVwqxmMKNhZx1aDrLXmD3VdvgYub3ZInUwbYlj6TLST+LcHKZiRv+2DsdGtX70RD1xnmOuFx4s
ZARlqkJtoPh8C6PVOxantkUQJMKDxQUXdDgcRREK83tu+llr8iLVXu1/bdmuj0ZPHM3DG8opz0xO
36x7/nW8dorm2gwNWhJnesdZEzGFAEBPuw/5Lja4S+Z8kWMstIligtve8HfOtp3CzOJa30a03OZa
FeTKRdNwp61BBTZeYn/mDu4QX0PXUiJ6C6NGoSjK5vVoSr0L2OvGXE9X3aleaQBmTpL5+HYzzzL2
KV+gMJVNdrt1+tbFv9PXNnPp+04OjA6RYTVcfm5w4Ua6pfYuRZKolfcVVypUbKS6uNxEof0nrpsW
710sZm6UWh6BPzbFN1pjoz8C2ZdWlvT4Al8A4t0wbt8BtwHqfDwP7WmdZh0OwI5nxtnzCPq1/Rfy
YpjloUIluUIkRCm6PdBtTZmFJCJ4ErkglBP9EWjXRPufnjgpfmLDzht5cfZX4UQ9nJnOy4Akz8pR
onn6OBwBqSnSOkPBZc9u4M70N1QftgJVXW1+XqgarchjQBgJc/DlQOe3DmFm+czP150BuZ/tBG5W
e0L3mYs3v4AhzmQK9nDc4X9AQvqC3X2l5ncay0wvQpQgcmBQZ4JkNk6ibEVxXXQ1vEUl+W37+gFJ
4mwAC/203x2gJtGrX36gTZvl4uXlX+h5cftwukiT5nCxnNFGXa8jxA5cGUDJuGfjSIvFYMi+7AuA
yjQcOBg4e4nqzYJx8hTODY0RaZdaFpxslRW7qC40GMjjLZLGZBbWG3kb6xuW8H6hj9wkyt5f9zkj
zPJtTWvesQL4x13nT0IvY1KaW3IyKt0r11AXR2u8ipB0JJ7S9Turg4J5fdUqOttpKOWtcNOteezS
jx/aUd7Pw+iM9V9dwxp1sGgbkvEaoxmpchCoa2AQwYhVyzR+K2lYjoZahrJydyvv7ftrioSoa+Fo
Wq7oqPKMAc1dsJoUob33yYY77gnKlT82lI+et1FvpzNRPf9WN6Ijlzy7LiFRUaXjxCuet9lADH0x
Z6BtL+DiFWMGudHQ5IlWhdPLdKulkJU+QWMKKKXiV/pZKdsEn+8tt04ORDCZsqYHjOKZ6uptPHMq
zfL1Vh3K8JiMrAOyzglzCqi9LdwFWVF26xsQ3kCefFGCc6NZyPlNnvq0qSrOgqBTRBu1vfo900/Z
myAWvumHs+ndtl+SatxRRCiBf5kwqkCZvNztr21FhqTOnsY7sLiEgjRN3432bC3f/8KtP5nmXDS8
Lzoy+E6sxVmwFX8vGjb2cDgV2E3kLcjJUhNdDmzi0SSRPAJkxBx8E2f8BdME0giIZdh7H8zCmq6x
RltXUzjP0fRRzr4F8qxZK/VL8fLgDb3xM4LaPtPDONvqTHFqeQ0CSLzfLCNRLk7QDSpHBJOCs+4J
HZJMGh08DjWGxJ5k0Di5hBK8WtIuBWNDe4TLWJGrryPi8HAO9xSsQQtE2advuV+HBX3DGEkQh5OA
FmLsduCyxKIxH3OddUFehDQ9LQV54mSPVv9nULFCVhRXlRDdWCVAsyMvFW5L6gBVQySYp4i3subo
OXp6yV6btOxaZ+H3A4vjzExfBc/R0Hz2OG5bfQK9ueamLrUMwdWV1+et/397cfxRPuKHaFz7o9wL
lK71tqyUWANzKJ+NcvaVrvYE83phcBHKmDHPjmzbrIDGeHtFYmLs9kfjglCyPAGy10iDXoKmGFtS
Y2hmwOMTIuXt7rzM7ZyO7KKZ7exHyOcKTRB7JGODYQmMNwTiiBT5R1fdxDU/HFfDZQ+gvyI3kPsR
c/jybesynoOSAusXIak4N3C0qxI2o8JLuoJtgxgkBCsSKAYg8fyVECIX5Ch8qcXdAHncVZELqtab
ZD8yCjlc6qdzPJorfutvumkn2dJFT1LC9uQcRabLN2SozxZsvYSuXCRZUQD7eFj/IosflYLPzF85
gr+r+Ue+LQrp2BCoCmODZ4qb5UG6uyq4uIIwPGG1W95wa//EtPf6Rm9RwTx/5HYug07JbP0vO9Hb
q6q/NTW7Swz4VktxoR78ZpG0V7LAoalHE+3QEE4Bneh5XsG59GtJ4qbbJu7r4xEIPQiN+3K23m4m
LzqQGHsqsGcZ7CnBdb1DqViMn0vXab8geT7pQz7qkvMUz51YM6ariBgaKMvkDfKbyw2+LIWBnFxk
FIfFYnY9PmORnDqdfIGpzrdcMQFM8AAT0zU6ZYlf280Mrto+7yP4WIX3RUH0m1Ra5pLxnkHqRlZc
CvVYqnpChfOsuaT/xJKs+ozhE+SHACaCKr+LInT9Dk9oSVFMLEvhhGch0YbeqkXP1/PNAtsDGQFV
P35s6asOtH7Lw14xacN10ToNu1PzYpgTnsUtK8vXYReW8lLo0fYosbAFivHCydWlfTizSjaB/s0y
b+INGvXozsKgUmULZIpqL8XS1blfAQM2J7cO86kDQvyW0f4KODLX0vVKRfbnkb5IB2UqswdacPjC
WOfL1Y+yxKrGR5KwIhM8sCDPUukqDrutErkdfapnxq/X/i/Qwa/hN1KzYGNbOw0d4NxQUClRQ9Wl
KUXL17yQKLeOic/btKtH6a0KSSiL4Cv3guCLNtLNtAxdvqR8f/1lJpEiEQo0RDbYf0/L6FL6/Os6
40koUBRUweDezhwK/3tVYALawURFrs1fD1AUr4haKM6ee+9Q8QeIidhTKZBWh6J7Jmk3VSMaRjw5
18brXHtLC3BVJ0oT5PtsqW8JxunSzz4zJbR7C7l4Qy93+M7Wtsm89SpyaQ7vTtRvo6hmh97E/nBe
fdy3cCi1r79hI79uSWs9rGYkiSIIxRvvk7KTB20HB+gq4ZMp+KCGwY2GpMlDGUaFGr+JqAWNEZBP
X8MijD5EYQIqfgcI2zoYe93dYglZhO7482JVsyqsIwFx2y6K38ho/kq8e4dJ42um8K7zciYa5h+F
yeTHGMrtV20xJRIpV/qPU/l5MXGJygdjzZDYhhKk/PB8wKvF2HIlg9pSKMNjZ1Rf+/7xH+0f4EYr
xR8fDGs1u2YFSrrn7PnF0OnHYnzthD45cWvEF87yIrRzJWMPYuL1Oa4CIFHxm0hZfYpKHgDoy2b1
E4IAAQlF/ktfYT44WaND4lnwqW48+r1uKl4zEZhB9qKl5LGujU2VruzWnKSX0Y0l3RJwZEbWiK/t
NrHzXcwbUyTInMkZWtMnIefXKi67ZFT0R8O+grPVMavhF46YzPB0QjvpAGMWzvnw4Czq44RDkhXS
WMfZ9jiHoV3nyF+JrTQdQbJwy8W1jfColsbau2XWpxisqYt3QU2dV+jmP7FjSpr8EP0YsRdx7hiA
ypYsP0vH9ulfR78zprBsXTazshCLNnSvHx4wXXDN0EYt9qIsdqdvuhyGHG7jhjEtuLkn5IVOMY1T
epyRvV13mDaMpBaLIis4S2W+jnbqbMs6uH03wKlYtrPTiEIl56/3OwCLDfLGyMLNXZBgCRaDW1aa
2tOwVpHDtfLXMGqWq5UVh0Bj2j8p2ZmNc9RehIx1U6ivaK5EzN73QESUPX98yqmTXzfehx3isrBd
soMJHjXfUKzc1xBe1sAnLtSea4EZd+Fb5jOSsSC3ubjyvEyT+e7H42vSs4nsZCbMsKKnGOi1Rn0e
BjK0qPC0YXK/1IN21wehUL35RQtgzSi2XYCnkaW3xue5gH4QQ7+m1KdQ2a+L7dadgZzWwwmCW4Qk
GnZHIhmrDffJqxpG6bh58/3fLzcf1i0KbViatMr/ehz79UbZTtthJZNxkSxZ8TO+0fpuv2dubabn
HY1SrA5a4cVIY/byXTOT0ZzykfD3EQFGfk2KMgvD6NAFEoPFuAb+XhEHi66+kUziN1IabT4w5qtL
7B7EwWfXlfAPFyGRF/pFA6Vw+MWhKkrIS2bYF1dfwlR0hTGDESta8KX8Ek96Jrr8S4Er65XxVjAy
je56LWZL01yhbOV9H6veCneMbTUwzBTKynRBL/uwiCf8Ci7/Txr5vw/r7ZkeUL/nBDd1mIVhaeoT
UOQN8RmwvsZD/6SdgQXeSua8lEdHHqLeG25YjdpMFFXHKawjJJ2qcvXzDRP8B/gRaSYPGnj917lC
Z47YqMZ8dmLcPcHiE4DVEkbcTL6jUgZduEQEZ7+0IN83SWH0XSi7IqsMTVKG++DG97yU35ifljPg
lz2Cnpsn1e0N+NubBlc8Pe4kt/s93UXsmpR1wHlzfOvBVL33R0erbXwXTpIIOKJWZ7CgDnV4Agbr
yZ5iRIibMCbbJQSmp5/igyOZVmURMkv7GIhj4ffe6C/itmGKoIWIJBUv6oAwnW4gMSNvfb99QeE5
MriJTSBii7fv2n3c1BKnm3L6iF10EOT/T3sdSTmRl4f0B6CWeT/ja4bak+z83wIc1T040eky8IpZ
w1M1itnXiebBvAbQc3Z0ibjrvlTq1nr+tEYaxIongIJV4m8Nw8xVf+MeGr+jaVLyvWBXVo88qiW5
CRH1znaHifiQJGJbGDGIICtlVhU/Kxs6fv3amPj8nV0pu0EYB2iSgQpdALlgMxq2gTn/GtoTR3nE
6qsdaNISWYmQVgaTXTkhREiVQ1V/xJ1O3Vqc6d05TPihlPBO3VePv7b9mjj494Jqr/ozPm5KrpXJ
+rmitIHMYPex6DW2l+a0gxash3OUiRXfhtz0Aci8tfYIHShM6PXUqb5yTDGvAzmsWKpJv4alpmJS
QW1NCb1GqifhsYSXosm5GejL3C970f06wah0u7//fUvAsZ3jXiTeDNxz7n7c8QwV4O5zqGz81To1
X6Qx+rzN7gDUyB5qjEiauU4Nv3TwK76S+ncxkPBAiY3lejW68yP+kO9LTScKf9lRbcLBlZrKMZ9Y
TiDx5+8Sb4n68f+JhDpTJ7KS3jP0/lyBtFtcY0KOeceAbCg0n7vS/SMaDauUH94TC+x0axR1lhhT
AJBwhQtjqoSbFkbeh8UfHWmHNySdqajm5YYeyQR257RKYq6V8g+muDHLOb+b67fai6HtOAbrflxn
aEfLD2SlhvUmE/pvw7NDBCe0qaluuvFt+YO9geqbojtke9iG3fsm8o5FDYEkMVXeiwtDANj5HKik
ovb/CtjFRkrvR+KS4L6Lv9oIAK6t5Io7w/prd58xhoghQPebQtMeYdmn19OztwFBVp6UlAZ7TLQ5
EoZ2FKFtnzXNZiSOJSU47IHDEUPYdjOH6FRIpYiENppHRcaGIHuNcySoRIJ2ApSLYfCVtMYI7om0
COfeXzbycXO1KjGyg9Jy2xZ05N4JLUI9PYIOc5EA2a9t2vG2AGSXrrfyPkGjO8r2MdZQCmKdKSmF
6R11yN4/UurkST/lELFbhsbady77cSAOMPneDBSqhGnmTFPCcjfI5X9QJYaDO/AsZygXWYJEKmjY
alEIQzcGmsJXa8WXuKR44kVwiBEog/vYg7zYBbQFdSLwKEvb11pCQ3Aghn9mhGb6KT5kWiICQlf+
p7op8a69goiySlw9k4mnVyTCuwlDFUuUVvY6UZsiVM8EbAD0Ime+WmU/hN4u4ty8FoRjG+ERXSG+
MmdtEBPOmqTl7TRF1iRJVEjGA2/kNvQbP7cb0nHgF1cxmyPNRNRaUABZcNOtMN3gw5vBhzgKQiIE
bFWrV7iUCvsSbEga8faMGPURcDI2V1VWMsv6ooVB5RDoAxE1WH5Iy3avgD3JVo/hki1CiC9R5Wqg
YDLv0QnjAXs0nnruSMD7lj/c84afJH/S1zudrNs7vQ4JbUOg1ssPo4lNrPUSHTr7wCmT+yp5MGCE
N3SSz1fVm0GE6jD/OEM2UHJx4L8MMS8fIBPi03N0NwC7sTp+kYz2g0F4VMttIyqWCvpPBkhU8id9
lA0aXJUYWMlQHpxkNdUFXFExxJip2aIdtt1vWK6pWdcKRL0RqMt45wwk6A84yjJiH6P9R3/Q/Eqp
HW3pi7GHkcp7mQqONgfv4Y+UhLAmJX0Uc4Wv1vIGhrZ/WHbTSi9JNEZugzRQtJA1cWmqmdyqAf1K
6/CsljmxZnG/9L7ssUZ7/YVbBX8CKr9wTm+h94q9m41i8+fmSJySyB0StYTh/IK8yELbpJpZwBDW
w6ghCpnWZJYDKsLAc+4cOdYRLoc0g/QICJo5kjVwwpyzQqbA+S7aNEcXM+ZD+dl5E9eXqBtPTVuC
LJQVy40hlLtTsSp1+WoX9HKl+3WOGSD1Zm4kameWfyiVJ+PZyt12njdqfExeN+JWwSN+3b4lO58I
H0O66W3Rb3A6S1Hvj0G7xbplGjfp0P2i2jZx/q3S3Vn++uoRX6iZjICbhArJKpuHQ5rE1vBh61AE
hoOxa/JN/R+FvBiejgl/Irvy0gNrkv0gDTEgOrwjl3VoLlfqZddZQrTRmzJLIXDnos44O3mK4e9W
4pamhh2UZAQg+0ocAzd6eEuUknTw6EVolNVG8IzH1YXB9TdHmXytQ8POn8S7C9NgXx6t/S5PQrhJ
IkRRgaFsmYLveAZqIwAQp0pvP2BzXfj/0n49WC6VRkFDdniE/L2VGPuwCz0Q5Whu5AwL01i/4dDn
JWWP0WECpND88rv4O1xOnZEbF38oTZEol1z8Iqstz07Z5f3TzCyfq1wfd03wE8YYz8VC2QtvaeI0
yQjHNh/19Uz0ycRWtvfVc9ggBO0vKWa4PptGwPlyfororpnQ6kqSPC9OA5+ONy9279AEr9NLiSmI
bB3OacS2v6wUDh8b2iI0RtzgHyr3GhnbAMOxjmPcGAU55a6I5tiTMRrpCNYmOietbq4j4/+n7fjl
x6HtzAV2seIIJ731ySRzRPiY0rPJauDXLu3HatWYM5e51mVW3d8+9nFFFlTUsWfvdjkAFVPdQtZW
86Hy9ibhBIpBBV4BMB5EFWJr+/pPNCPKnqxrQw+eDQS/i0jFGWEAlbpKNug/9U7bHNq1umqtFFIS
pJ8W/dFUDCjU2mCZbiaJmx/bIVKlfh7qOacioP72bC0yIyrZro79JJ8oeX/spppmtOgLXWeQoeqG
gCRuDPOibtVtvBslYqsiDKWBwYk2w8+SpS/SccyiZK1Yai2pdw5bBAYk55PVKKAmasu620ojjAVO
K3N4Q/UvwQEqcLQ60Ao2EBoxDEfyi0vCi2nWQpzLpFYw2aTK2S7woOafYh8BTxsI331Km/mNZpTO
CWuOIybXmNyqpKZLGgGaAcxvE5gyJQCDc6Q4MOybR8KluOOD8WPM0+t+NFQF6fflvlFSGXfDn4OO
LDRrJE5y1doooVWqmAIwGZJQJAniWqh91wnsofh7049hUgaM+z59PjK4oUZZfsrzpejMiGOTeyPb
kuwydpmZoPBws+eGYQmOfK4+5nU73NP6pWtB9Sk5qbNbZ6rObrOCo1+HCT9jgtQMEXdGFal+Xtd2
wv29mtnwatdAPIu9Wxwzu7ZA/aPxctj6rCUbX2rGO4RcIoRZiXgTzDip1z0etTRKeexTRSFrG3Hh
LeJeETqci3f7X9o5L0LZ1ryNq+T+GPQGBQv8XgPXeweRIisWqMim7XW7euwAzoc+oxnHokqIUAO6
3Vl/aJYWaXCWzgDXV7ByzWl9ST4uLL2G6BAHc3jqidhtBZUye+v09C5NUWIiwemm2ovLubs2hmJs
k3txqHKLB0rjlagYrtqufyxpZTz00cP/CbBJklrt5ewJVY9moyT2Ry8SLEmLn/I9nxGgVK+mtzue
Watntj/zl4zoM3jv4caXHm76gdQ4A8yrNMglRW9FMt4cr6hN802d2tHdJnDkDO3nqsijjr8re0vm
P93KkgQ0ZMrdBUBiPg4YuHBEAB0btF7pbxyJ3zCjxb4gzJ+yDxdHYlBzRVUX66X990szdX20JNRU
zXCbnGV3w0d/hk7886DtchbnDje62Fcobias3dm31KuwCi22hUoQnZGxa5fskRrqDZjIsqKhHiDp
PVN58Ex8EwCi7pk+gqW1fod1clTGgRXPL0+tHF23IkoBAA5lQIpbOKuxKwiJprTaMCd/LwZBK1Wr
rqyqKqlfBSCkMls3JB0zOAcJ4+2xUnnZxuY17juCX2xCHb5jFd4zXtfFIDC/D9axXv5qlx6pUDNc
GY9EkFqJu5flzYDc/XleTkY65WmkHM4u7IZyKZJy8x8owuosJZVgJ9G1ieHhFJzriIEmlkYIK5VQ
3Lofm8GXRC1vfZhe44qKj3oLgzq3zOAZc/+Ip4HzIgvWsnKM0xHvraTIxDtQji8nCtenR6p0s4ZB
Cs7WZLXraJG5jN/X5Vgoef4L2MpslBkrB7pGPognVeq4/sBruey7sxMB7YWvp9yQOrfHNq2sdrdq
/fV6ABtJqg7shJtFyLPueKGxLzntJJGS8RL0smhgj7JqXubyrMYoOeZacpcTMU9DryMtvAexU7hT
JPD4OFQmaRdx8NdYZkIiPYPEH5cLTKQ+uwUJ0znLN8IlfVXiBs2fZCsYuUOhPdEqj1r5AT5cTDyS
+YZb0PQbnWhiXw++AEO8Zc3dHJL3JIZ9gtqXaRghH3KLEM3xVSO+okjaZs/tBz6JucbJusbH0uHu
NGixgxEiVnCwb56EyoxGmLpjVeX1JWg+wYSozm+0KaDUgRGVcUZkytHAYpcFOb9UKboh24ldvmFT
ICyDNDuNppgNU0hxoWGTy56t0dFVD0VFtZ4KoLEMewMvkQJQ4EwU0zEhXrkFr2ucI5YSxgUwRfLr
fRae+DNDeemWRnRDyaqg6wRjCEOUwC1Bj7eZePJGGh/Ssr795Pm0yY8wTV8nVTnNJsRleBOkGuu/
Q8PNzSTS4vOWn02aEe1L1WF503NMhosMVbdNJ8rMb53XBtwSvuQisQCwUFv03n0MjqDzQZD7YzSg
rsVra2VO7vEdCQIo6emB7J1sqJVskkXnsKiwka4pztF6XpVVUIQGBeIEqvGR6/RvXN/lbsqLjPWG
JAeMlJATOoTx9ZHCgs9a94quLLNXl9NJdAF7MjQqCpO2sp9yHw5VQckZYAC7r6Z5FJLKU32aGfcg
I2Abi6CEjkvv6zu82oJED/GWPiy4Oxt1/BwZTYI7ZpORI8Aei/G1Cf8HBLGN+inMl3W8MmKjnxfG
x4ku88abf9Fp4I9Z5B63snD1HHS6y7m+AR+iGrRK5/6JxylBlXZzWeD/eikpv0fC7kXOHDBmdqmQ
7cCSov9Y18blJJomco/8YCJGBZxss2bH+gWod/r1qxlPpqXhANVyhLy0nAk88DVkPRy/Qp6n8X+y
HSdpCq84PKOWG1zfXEFKUUNwxSUMC+Ek8lj8ZdaKupMNDcWGd8A956GO/7eKbtvtKQEdLHv67rrH
23/uOYGGWkjpKonmN5a6z33ogS4E6wEtkDZdv46bU4Cd63Wh4Fkdac/KStiARDaRUb5rbtHl2gM4
AxDoVqxsRE5/BEAznnlSGQPBonBvpTMpAcBmnd2T9vyJ+Xb6tzq4TqMRK7x5X1JU2Nfotn5L5N6P
XwqXa+Vc34HDlwfv/BShND/DhxGUxgHIxg7KjS1YRQSs0Oa/JzHg5mMd3Qg1OmwBSsBJfoJhTdQl
o6kKg0B9yaq/vMlL3HuL4Im+6W+AIA2fnetRw9iiHMPC/9dRJLzGHE8tJv3qIAAWdUriTRPHJDA4
H2qXj+dcrRcla1UhJTtU1e1/5lRNjdR0qyMT+41r9/xrG82MtgCs7X7SbrJkMP2+z7J5ApCCadRL
ZXrWKSSrzGwidu86lCJugn/dE1gO9rotxnf8I6xWycywM/ZkM1E6HSwnhK89f87st004woN90Vbm
nX/9Okfz6R2jnnKQLfYJsjuJhkK2FkVROcHEKRU5mHCPWxwvUVnaMbh3K/0hCQhUiCj4mCUjUBlQ
2rtyxCuGI8ITSrcvRpSKuRlU4VEmkagMvjQzMx2+BUR1fpvjCdAdcKhg3pnvLk1Z17SgiVH3OMgd
ABMRRfCaQ/Ms02A+hAWLFA10pzyqmE4Xc10W40ZL6jOsxxf2SNE/QRTfT9nPCCSCwo1kseczs9En
c3pVXILE54mOh373Y3UO18CNhEatPzP3wOQX55Dt0xdTTnH8vd+AA3pqJOXUzDwdkipuDAT9vtpU
3owUdG5qBMfoSNWQuw7pFXtnuY7m6BRA4C1GALw3hx4gv9lafp/XDBLXwu5OK4tL3geTqPJEh/tG
oBM+hiN6usY60SdeRF7OkAf7ztqOQ+WCp64JJJdEbEfoITy9LIS7dhDvlfvhUaH2HmmUu7pBsfY5
Uk3FaP+0hXMuOEpTlzSEJ7GVBfF6yEwHoyMGfPJGJWBMjRPk383f6q7rCH89XL9Dc7kmlwB3Dx0z
kr63eOGknCyCkY7V7vAhUgTiJl0iFiHeXUPTet1z884b2wzwAH9wiMgC6UxayrGQPoLHADs/8zK2
zOIJI2oAO79tgIVoyiBD75mXhXvxljDMF0AkT/0HxdsgJJy6L8dyJaYp6/Gfm9VYvbbsllsiflZL
acrKTToL/SRTCsVSxDz+i0O/lhthNdpkVHW/ZZIlG7Wa65B2IVGZaIfgt01zy1tdwSRMjtjphAas
XmN8fWwEWRTtZEyuLuvlgRv8eTzfFuJkxwArYk90IsoHDaeN63oKafSJQhIyQYXAG+jmY/mZB++5
uhDFXR4ereJGoAEpFjgOsxajBTCEQfeTvAmIlSf8BnrEVWlJoT0EtrmTv0BFIIw5m2RiQpVLFRIJ
w3tZMfuG/P7Icb707+4AMImDw67NYf6t2ysDDVAkdZWezL2aZQdwweS4e2qfFAqC1hs8+n7Z7PCF
9fmiY3/xyK+py2fcwaPsMYaRE6SELw43pJnpvkXmB49DVjdmZIx4IXPvZmTq1X6SbFdI3/drjDe9
ZFJBcq5iCByWPFclDqsrwEsnnwCF3wxDYke9njo+mLO5CbCmT6Do6dypyH2K2Up35AETWywqZ1ug
pOFXAGz78gJlpC/IHr+ulo7Yp1zy1c4bQuebKrGQ9nrJNvuKm1fZlJzqk7OtwD3rx9eIAKnBbWu+
RU/MBb4suzpBtPEQV7e3Z0nvbIMYaCNK7ESPnNYo3Q2ecmCayrgOjMfnL0feCOM2oLvimZS21xYm
niL/CTJqEvoubseY+nuCu6y9jGGojP6a8qSRVpzi2OkL6fPH2W+i+L2ueCEr/zMoEekIiHvB8Nf2
sa+Qo742wcinA8qO1PjZGbvm8OVDRn8NlhKLWHYx2CKcQzON0uurejxCz04s7UqchRwjxHW3K7r+
B1XcpVBlD/ILw2b4FuhdIaO4D61N0bJeuNGdRFgZCr0GXg/b21iQLGqR94hyvn2TjIp949G2SNaN
2cJNBcQRfkmZxhFUDQbS/ov04KiN2mTdBMp+/sE8INadOSHs0CT+YOpK0KS+/qmp63bkm4IN6VaJ
yqsBR2xjTWRfw0l+0efIIBz5dt3OWVd95ieAAmn8bXCT2CubX68ZvSVzE7RxGhpOSY/o+sDfZj6W
Fw/wGxNvcPWdjUy5Qu4dh+6STutFIM+EMz3kzxMGl+Fxepw9spMgu8Ffv6YmWfi/8csv6mPtrFXp
cncvGonuQ49YWz5cR7pl2foVMfYgasKwGGl7RhvfJrjp1TppxkdSgx4AZX58xgwUlsK5exXkwqJE
j/6qEf6IbztsFzSpSrIk9iBSpEZsPJ/M22KhtIcnY2f1QyfxlyCCw4XPWLySa4bxQb3hIKm1rM3B
LVMywLLfMkYpEr3Ec9UOhkWkAtT6ggtkYgUjh6I740wO/+ok20gVbmWo/Qu85Cs8HIB3ox9EkFJ0
dJChaY4K3YQiYKZX1+LvgMuyyW4REWDXSfuKZ3+ZtdFvjyoBnVTWpE24TpkycFb24ysxS+4oEq9A
+8f9u0SJygb4O2pTWH6u2ohc3C6N9sVuyCQJeGngkaxZpQguKazAD4u0/y08K6L8E6ugD8zNacq6
oNbrBYe104b/SkgQcp98elYWnWHfl4n/wEKJE2yg6fwM8pMUIIOB9Jhen6DTjadRKKgEj6eDZAqT
g0AY75GnjOwg2W+5O89JOikY427Bd5gq/OjM+3/vL1o2SHw9sMm0LqcjTliUJztCnK4bbkP7jTTo
gkUKLn5IZ9u08BzehBrzkdMZLxgUqIHA4ghvI7PrNWVtZ42tDfR69SefgFQwPYiG1eaxE6UFO1fA
mpFmqdvOi1+4oCu8Vs8dLB1gcPM1AZLUlXLC5Z9cH17CMXuUmI/IfOVnj3jXHV5vQA4OS5PMDxEg
KIxAv6vGOUIL1/zzJU7rjUvoYoeAxyhfGii/oChSpMR410soI/NvA43y4VoqAz7sgCnt4bg5GyhQ
HRa97m0H/X1romWzex8KM+2rC/SC7I9h/DKB+ZerZgMYAqK4QgS13GDrevCmHBinBuuSh+VPPJgJ
rnluT/ln+rIs0NKSQK8nMeAN3VaLBOvXbBB3E1pKneUjYGQDm/2pwJfGQUZML4ximafOdcf1uZ2q
AKBuvznZ/IvQkD7PeTd87/HT9ZWseRVTHtRdZ4mrsu7PqAlFoKxCtds7QycjLllHr7eRCC9ajRRe
93unIIT9RyOslD7GqeDSvChmMjyrQT1p34YQlCaEO46sZXhin3Nd7xwJ1GOFZneQsIT+GNwspHbC
f0OZr3kZosUdyC/H841M4+HP1YsEwEo3D9VYK56t+DQWtJCapZmJ+WYR5KvNwOWwbko2YVVSJ0mA
aGcQeeSg1Ae6/L8m3tJt2aFcONk04Y2sZE2A4m8iU8YFu3tpd46jf9mCW2NIwmz+2f5mkw037uJj
Hh9aKvSyZiEJsiCdZSSH4W4/F5LBWjt+P9qUOPqvT23CzMYQJOBty4BHirtfih7Npv+P0JUxSs9l
+EbPJt5DdA3t7EiXDud/1lxQYQs7pKcl750Z1FNFixfoTQSZ5Jq80rjIT/mdnaR+goM4zyvOLx5H
YtkPtS64tIWFPXZYXtnohZiA4lNqWd+pMJvbChQWpzRGRcDDjOUBW9CQmI79FghjgoKoP5QBQOU8
ebf3LOlQ45JxXLeMdCYHnSeSGgPO1IBR70KLXvf4hdKqAT80aNS2WdH+e2CBhhmur5eDoRfXeXiQ
jILZhaTWVonjTNmWxVAKm9Cp20DfLwJHj7WfUO1sjfkXJJbuwHqSVm0w21wxNNBb1fuebbu3XhqE
LFy2IyDysl4Mk+2M0mTuW3dJPm8j+U5suSh4pUyfiiBdN236lww/9w+b8lgfxBtw0zjfeW+Cd8BC
suTenOf2f7WXaBc2vpUORt4cOnek0bdA/EyCcnNC9YHB4goehTpKRG/3qI9irwiGFnlY8PRlRMLG
TJtNdjS2WzS8vv7OP2LO8Xyl1qmwy0OvdwNdS9S9rcbMPTC1wLIdv4htSmskEMf8pjE1ak7Dfj2X
TNWPrmznpYEtCthSVmblBBbp4NO2eOmXRgXJS4hjBBl/U7SYGv3uRgI72VOe5c6jfCjtngPkVDUA
zSnxzudp20MIWm/KdvWduYMRlIgLaVVgCHp+S2Dkg7iPMD7oAoDe9Hdx8anNEGIMKm+nV2m1dVtE
/U1vGipt7Q+1w4Wdsfr3/AVu8TRCjYoqrmX6EU/3qfoHxp3W+1SLS8MQPpVP66Ocpv1X0Nez+XSX
h632yv88Vllnubg3ucqI6i5lJoy8dp3tlJqR8c8rVKZhXOMWk4DyacedaBFZAi2MYRJW4eudMGIe
cvU0vCZYbawW7bC8xLvcix4KnyBppqTltC8C0Q1h5WWBjcZEIbhCufK5OPjrZsgGYUnRoTHktaBu
2Q3mNiSYXp1Nbfkba/d7XrDVi6HwTY/TAuZlf7RgcM1cv124/Ck5O7AktmktrTfvDdWzBI4kriAS
FQlqvJulvPD7vOJENuLN8ii9tsheomMcxkaT5HpvDtcxgl8GjHu8FOitHyQ0d6TKOXABhE+OjUx1
XBZVmAUZa5uavqpJsRrLn+GEDWdvVtYWAfAy9eKjIViTOX5OnYrTqLO8xyilLP8FjSx24jY88tVo
O0luI5Olf9vq/Vy68ChtM3apvU7jmoHn2LuwZM/DNR4NhpFImFAT9sIC+M2gFhZdVSumDkw8xxXq
srwmmhPsgPeLP56+sYRaIKVPLSBYwJjipC9pE7ig7+ED/F9aLV5kpnjxNQvM7Au/2a7bzbW25TjE
y5jf+eELy9NvC+4ak9lIgsc8s43BWEPFQk8Jh4l3C90XVOKfIc4rDpulDbv9tjIS96SH12v+wzeV
whGalilHFxJRGqV0y8M2kdjo0JhRk+PI9EknRu661eVu3lpwHqTjlMfqtPTDpN7VNlSwGBpzjRqe
nkjRNgu0RKFPesCLzSA4XFsKHiBuL0T/GX3Da9vm6wT4gkYKnPPKTciWkoEGwVmxhprwWui75Gfa
ALBSh7G7g3NGHf7Bm9yqjlxld2xCPQLL/lG9Eua2r3EzRxlR1O5UCT+3qi9iqwNOwcE/Ltp2hN0h
I3MVuu61DacH1JktpybdsS50Jkenp4gH2q52nFLc0zzckjbBicTdOSbjT3NWDilCo9oTCiQQdLpV
YQDCwTOdeuKsuA75uOFrG2+x8peWeDec+d11PyTFgXbFJyYYCyx6SUwbI9YcziROxSoxuNLwMXZ3
xReDo7yja5OcrohZaY2IRMOAPlg88UsdGj3PYn7A0sUCxdSkuQHvDdqkztD1iOHE9qvioldWoHM+
7SXQiZW7WHAEf9oPcf0Zl6zI/WEBirU2OcmPg9Yr5w9+Oy0KmRCdRXqoIGmutEIx5uK/Hs7zAM7b
0NiTBi0V7d+DyhxVjso8SrBXCpBw3Iu8r9AHywB1Oj6CbmbWWdBMoiGQ1TYM0Cklt0bEgPgfHumd
+/+/VS0SuiWRrjpXspbMwiLmaoHNZxZ1do+T9QwENDYmN6Vf8/uFZsBH0GJ5B9sZJoha9rU65EwA
6kXX/ZxJ4+fIv+/jbdMaxUqDJr6Ou/hmgcSicwZVFQu81GGlVCYp4HppmAkbJkHs12VdWbgJu5Pu
ezFFCGKPiKdVYzwhGgF2bjq9qGB0Iyfk1l2i2FGGH/kYSwI8zX+z4Sc1oegfVDIYk708wi1jztdJ
9DQVD+sSwkIdkDrXfXkQX3Wf7mThCKlKLZahY6zbQa+4qVycsNkES7jm0/9272oDL97JRkRBgCpe
koHXHOpvCjDOpAnEnY/CdUGNI52sLSnhD95GeKgdu4VT8FFRMTbq8xQPor2BT/ZT7yCSnaqk2BlG
cOfVGheauATonDjmhjEk/UFMCZEyOFMVWvs74Mjh3RM8O6bnXLFRiYa0jmjMXeRPlQ50WMfZPYeb
r8zGq3QYJTswNfSJ6FQ6WquF3aoO+FJ8E8Q5CeA0BRgqy0oBKTyCxnsvips4lwWrEzYLJa2qMiL8
jJ3iQ135+fR6ClMZkA6vPvM7On3eCBc3zvSm0+ZxxtclKsAT8d4AjkO3E3TcVqh3vxjlLJVX0VF1
JjrMbtitx+1KkrlFxfiTrI/3UCzkSvdMnkF6aNn0334l6qdek46VbdXGYrNjJzO6ctTTWx+dj01V
Bk0wOTsv+v1wfppQcNhVG2bv+HtKNdg0qA5AaNnA5nek+w1gP413nf6KZFoK2LeVkZN+ooDxJMKQ
RSw2/IIVhFLNAC5k1V8cH8JspYqEVyGsEEafYJiN9O4wUopLiGvCUZyApTubHEkl+btwJZozcS7q
IhsBs4X0B3v3XikLBYsK3VUXm3ro/jdkTp/vRjpbPAMoRaQ9Ln+DWsUOuAqkxcdSP5DeoS7m011o
uAEmW5vgNlgDXkAyYscumJO/9BEaT5YD/70cLlbYBru5FzSznYJqb4rRMUU9wdGqo9gQQeZhYpqO
pmr/t68Bafx9kvuz6B6HZptnYduhfeKaTvUgIRs8UMA9dZ6N2EyY2/FpCWiAN0k0kNgVlnNve0X/
AQdG9jt2HR3GGc+wCM6ywF4TgYPK/hYa1IhspFaOyLF6VDwcNho573Ox6SLavnpFJhqgcCmWitCr
U9QywBeZT70A4vF3AGeSMBEFRchvy7xeaHVRc+iBx0KoZCm4985E/rUmgCeD/8hWl3HSk9ylepo3
fce+kf56a2P0wyBeAMd7JppCEG5xc5B+Gdd3/7fqXxcUYnOghHw5tZonafwl9b+l/5OYAib61n3X
+wV6Y+36WfU0V3LJiVN1qFTuJwJHnU0DuURl8JIyczlHEHObW0B1peDHdC7yMPxoBjTPlMfi5HUM
mGT/9W5Q+MyWHoyywk9CjSijk4VFZCQVdYxem4RQhZJMtPBPmEwjM56nIXqEGsEDkoGw4mJOhaJ8
8wAg6obq54r12REYAK2fzeYCNlh2Mb59JLjYii64QT3W9KCVCqlk2HJDlWOVhCvu975+wsPp6HkJ
z/UTR3uWJf/4OFzquwcU80iLiYvkmVq0bR2M2yftzhkxzbm/G+BmpyrbpYXkVuYZpZpGFEUXuvdZ
LG5vwY7y59gG0qqTqsrpA5X3i8GS/UtYr8thJsFBjBe7rUHhPb0VHxrvAYtMSQX4771fwgJKBEoG
7AAmLOEvvnAnNN2v5rzRBLq1UM3ZNK+4b1b1sZe21d51EZbnWt6j90/tYXc+i4aR/zgQTrmejy3U
jmCut9PBphvpWPBlgoKySAfizZ9yPllh7fJb5JuXFpFh7QLPe72YtJDiZ2Vcxa/rzEgngmedAmMd
i3sO3gz2qY4pVT3wUeGJPd4zYSvpuA+UGM0kMz4aWAu2qQ7xV2RkitnmK5qr1iv8zgs0LQqUy8YZ
D9t4Qe0BZDgVBcnPfC+QaFhlDHHcAu+aznPzfJMErGyihEFLXf1fxct0CF/VZfzCiQJuX0Gta+zJ
dfEdj7JE3OeUDRy2bUF3uvmnlJlTpN9bX54tFZKyGSFJmuIacBjdul0vOqu9aQmipTQT5flJiv8Y
wM5Hiu8f0os1PjZhpe6h+26bofrZa9RrBmMsAlHHtFb8p9SNLPKRGVka0nlNb8uNWRuM6C2+n847
YC3knGw+IKavA+ltGoHJvyCaJSzxVJe7J0Z+jekjiPlKPQPEVTVA3t2IO9SndC00jKx51I4i+qu/
lVuQ44JtmOymu70HzcG9TFp6lJPJjquuWG4avZQgzYDf+i4ipB6grvzo6w4Umegz3XgscXPccLJa
KBDS6I3XwkIc6Pam6EdeyfL7e3QFDhft25xLz+p9KWf+VpwIug9fYRnELGzi7ukNfVJnmwewKu9g
G9D7WxcUorakAylfYsMcBscIa6HL/TYPSKf7CzTNrTH+HPt64zYvkj490WbNRFatrv6hsEN1kg/I
fGcPcgBHkbFfj3QcPOvIjcxrZoYWXvOAFtqJu53IxmWhAA/6E99PQ5qJbb4ByQasgliLbJbymjSV
4uJxd+NxzNpmt5m1Sl3TykTSg9Iyxtxr8I8n7T1Kz+A9dvYjJ5fo6pkwpqSGy115oXz4hH8tCpEC
1nSnnoush71VOzx+iFoKSz34e2UY3U5S1dYO0wT5PKAh3nIDZs9gL2aEKzHgMK3fxs+kFuvkEUT9
RcTFH6xp6hMqO7TX/ppAOP9udp2CG3sLFflNEdFi89zv15d24G0NYyPJ0ytTEOn2pPZU0Sf6596f
/QAtJbQYR7e11bJpaZL+yzxdJvAQbvtbU9AvMmsJbcUgmfeA/q5Id4sxpKVUdPWi12K+1Phf287G
j2F+Buc1Ms8giUi/iDSjf0xNwxlXoub9XnjnRDxa496++ztrOsA4A6cBs0DGzhYJLTupk15zZoi7
HNP0/0kO2yuUxtPI2NGarVr7womnct+8UYKySlyhuamiNKte4WvGdYEFZ9jcxlbm0Eu/qtOddvlM
ZgPm9H5lpzRbaU+EJl9ZwnK7vJSOpG0mIjHp9B7scJlMaN2RbJMjlkyStZqpCr9ga1g+0R09Yvoq
CsuKqbef/GVb2CsV4T8ChHT6gLR3cVnPvttl8muAImAegk3a0wm7ssM78JbZFCttJgW7RwlsrA2/
H1lv0t0zg0r35ewcMDi740XeWkN6UOGFkUFcbT+f1IK68qhkDNccRtdvB97EW2N61T2fUS6n8ZVa
NhkK+URav1dFd31TPgZPZWV4Di4VB+AH4+0ERTbgFBHWoMX9ZaxQulwTvAJHR2QCVrb5v/Pw1ukM
q90hbo47kcv2XOitPpTXicoo8j0DQzZwbS5vlT5Nbb4TkWOIKe242Nim9GnRCMDiwn2TpcaLn+KD
TsF04GoTJVqs3Z2VbX2ITk5hhLZexrgZEHpuOZpNu7Xcub+zE5ZOouE2V726Oi7SQL0vAzwfOfKL
gM1dEILKKhTwF+qu7gdg8YFiDGn05dSZBoHtzzAY0cDQRabnB4FaTLPqbiv4kFWPG0/Z4i43wsmY
+L3pvh92VavJiwKMnq3f6JJZ1lqqV1Q68v8kLAhh9nHLctZlWLWK2l0zCA+U4FNSsWaUtEoHZ8wW
pOGzXAGZ/cYnNlPiNinDrguRd/sXzhsD1Sx/2a744DMzWfZH8H1mMIqMDQKlhId1tY7/RkyTwd+h
K17FSd085AAr1xAUpNWp7z0SjliaZJ2aoRPfW1jGJdhzo/xwR8CWFMcAox4IlvdSkMgPPz1b68M8
xwtjTMUWPvPCplBFqv9cQ3y+J3MQov8fn9e9yzOLWGu9mpHjGYIZkjc13plExkxrmnxd/UY0vkwy
F8XuZKtYvvZcEo7VjEOvM8wa9UhlXh+Nfiw54KF6eQkVby1y/GzGZF6++wEkgNEffMHyohH3w2O0
kabJcL9oyhCo9R7O9rk0jWQ/bq3okE1j/OFoaj/WixNa8yL5201nCTgCMxbvjdLOWlxuX1y2Ea+n
f+YpzOz12bslgofrA2auRPnVSulqT65bOCILNy8c3kxyHrJdGaoPmihu7dghiHe6GiKsYSvz+cwn
NyyQ1a0bdD1B53E2WrTnjDdgqf9Q4zUOCwkN8ZlamRm26EbpLOzbUmytrlksANlSXBzAuiKvdLct
PGAKK3ybxTU/momxVXyaz7DubJYJk/xV6V8/RCzfWHhucYjG8YbvJAZLllj+NcBE77mDDwKEJ/mJ
UpJNs0rRIdFcBPwl0fSBqn+3Ke8ehTClgw/ru4LLX4K9ek+iX0HwTcYtGzuSMwvD5riSXKMqeQDf
jS7pXjlPWFYdehLs1alGUPC1Hyh5yuv1QF9u3p/eXw2Z+trx81t+N8HhVdnzk+KLURblWRK2LGSu
EjFv/up3vXb+rCD+YCJKc0Xrmx4bHUQlGjMkmBiraOS3o/QxJfKK7L0yBYU1DxLFwP4Ph6Y2btYD
d5idMV9qRMXvWfJ3CbSkSPWs1sDef1IjnaMgBvoLiIx5d+kcu6gKzZHjA4xnCHohyQSs35+jfuH6
CeS4Dd1e0XZHY7yPugL0tQSraMrrv/9wVn2GFRrNjVB3bGAMcXZeOZFjDiosxuf39cutTvNIn/VH
ErdEbowxB/ZWAqqTjQvg2b98OJ9bieAqNQwHzjT2T+mRqbT1k/Plwov5ZwAPF5YnXTsbUkc2JQyr
OHE+aT3aNQVBbaHcaMVnp/u8EapYdEJLKmQ9M48GxU2y8OBLpDGPxKAJZrbfbS8n0m/UK4ro/n/o
S/Y+jtrkG0HWTH9Jw2oTzi65zcM5BcJOuMgco5ti1b4nZz7zKIH/qfzrYd8Z4J4QJnQ4zJVUtPCM
MXetZXDVGlq/pzP1c7yYcdgp9O1Vm6tMfQoEpBpUMgQ/uDzfCNM3QBPSYH6xG+uCtCGhWk8YUMh9
5tWlpx9S+Vy16wgRlYRHmKlOtxsqDku5qXO9rXtwovkvzYbVAY8YndRo0YmdOb1ZGBNc4jTtYLSD
w5qfZOExzIsmMUzJsyfQPkCiBTdyoUJw28dryg4f9K7avpnR0nEJ8kQsASET+pAdEWu5izpBf5b8
USIYS2klyWwhZHGu9kFhbJ4tz/jThhszzJMFGwjsVXgAPN0pTifKtA4UmCdob+g3CQG9rGwppY1m
NZ8E9G88MhfDJQPf1yexNftGKiu6QSzYUzGlMtuM+i9u/SxfF5NUgPTCnPI4g8+AJbJlGN0UT1SJ
nnxqGQkr/z+PJQ47ZQD/pPZEsX33Qlz+Ly/ko89dBjTxnYK8pLt1NuZ3X/8Rru3o4lUaLQqsY1TD
bxsOfsQ7BbbtMaTemi6aYB6fHYkZ+NvGs2TL0BgrWUmWa8DxZYF9FTQcuvohu2OdK9f0CJJFlEzf
EnGDMYlfPdXESlpUHm+h5MG1UkeXf3K/j+NoBcJc4TgYZPidnjQ/3zJnnpxJmbfXyNc8NTsRPo9c
3lhVfwRsLN7pCsNwPz7qUnb3EXncFYYo3SQLstfcdexrWXFwLWQcd7idp1Z/BZCRKrSuxO2vzy0L
ZV83lhuCiCXSwV8KJT54JbiQlI2EfCWW+F9UlmPUj031PGF3uPiWSahvzoA2Khb5uCO+a5qMDrDD
dRmFTCUd+JrDE8eZwPUGcZZROvlAIoNB5CJAVGGKoR8lhF6iUF3zMY4DIRDpg7dTuYgjfwaBvrYs
mPL6P/cb4etBaG+xOSbki92l6tJKGPRRMgayC70eLVeI/Scnkqp30hwxy/eyrUL5Gqk6vlGh0hyq
4+AC/OuxTBmVbZ/xex+3ut1BvdWxN/bWQ6uKo+G1bASOae6cxwIF2AHR0lazZclMa34/4X2T6z0b
gwRZ6YXmKL6aXJKzbROYHy/PjSZGJH2TGp7QaTpgXW5ZwSFlBpiaLuEAO4WYG9dqCzoGqovmP+3A
rr2utZfhWFNmqyt9YHPrg13IemffxH9ikEkluMz0Hu48wwYW/d5XlnjZKeR/inER2zDiK6ajuPtm
QO5Uw6fK05mMw96hHg4SFGEgMpuVJXmHRB5ma07bBYpAOjarK4Tm56IBKI/aoOMxvGmXp3z5cQhP
BGTzj0Ih7V5D2USlPoYcfWmkvyo2BW4bD+qJDhgqn8adIhaRi59GkjOwP5P8ZVzyr1UkaVtQASy5
nPZ4ZbyUvYMqJbM1UfY2X0hcO94mGH6NjVIrptZOAJEtOFh+rFmpgv5QzeQTY+hTqEPxgM4s+QLW
DSv9XabPIHHBMRianInVvzpc38h6UMVh4iGkhouYu9MvkpOi0G/PPpOKxAwJIqrfurr+ab0KlMCu
2zd9942Jc5VWiJ7e0Vax9xkrocqy6kgtvM6QOXsQ/KFEYpBNJXmESr51KlmRq2S3uZ+xbzeahDma
Qyk1VCFBb7tAP5JLY5NWVUL1MdePxrNcpxjaXKlPKPForQu16bODjoRWOmZgPjTKABigErD8IdOP
kJWeL0FPWh+UMVublGnqFNB24Bcaoy+iYCUx64g5h4QOjuT4aVzPHIk2eaOhXcuAB8KSu7KTfHpc
vywGsdFd1C1EkUYubSdoRGO9y0zhlSeg/6YnL6tkxy7iQlkzWwr5sa6R8XN0YG8espGjzLQuXQPY
ikTcuQ5sgAjV1bSXikkANJzE8tSyc2RpbRnYIDnER6+to1dOdQgxck+K0E4tszvgDc7Z5M/X5laz
W4P5e0FLsAz91/ZiiIgaC0Yntv2MRNv8+JDuE/OZS4aJ7bbB2jDs4TamNYC4FC2Cyf2FNUh57rQP
7tl9TkULUNOoHemK1SmKJ5du7HY4/HeLWBdE++qtojvCznPn6GAleC7Bipj7i1cG9qCyiYcSggqA
qdm0tSddf6xElUyRFPbQd4uvW9qTZVbIhF/8stl6iV763gXhJQ8nreNeTNYgcj6kuSXQzrH1BKIQ
Bls2eAj6rSX1C4I0sAvfho6tlJ7RNhwPW8XvCNRzvJWK75HK/r1VXRiZZvHatG9WVM3St4Seb5hk
vzNMBj/iKN24JphP3mIFnGyjOhESWJxaq8DnNbLLM1B3OPx/57nIE9t8oV7S8xESzaTAL7UCMkXn
BkW9Gy9bNVPfN2pE+PNlMcKqtLQ9GDiVgqeys5q4Zkq+UGjwKpEAUvJIwUcT8xRh+QUAYYMfehVy
gDWYOkhj3DJUMOvFsgLO7FVepdGbkw45XR2g3QrPfOwOvkv70IOvXXEcEDXYnmq6ENreAZyAqr8T
LYV0xSLedVRBTp+q0qBmUG2E0diE1OedXwopgHtOM3KUiRFD2ONhIu8lsHv9x96U/B9YHnP9Hubf
qpKxHZv95vfHotvnBc0hCsYkPni1TPnHdH6zkQcCePF0/s6cIPAb3DHc0gpVeN381Pu4Fxyd942w
FMC1Cxnir7Db1XagvPOom7LqhdUIuKzh4IG0Dg7FSVQd9/wlSy8Ga9kSrp4OPTDrGOlwJzOynSIr
qerUZu9jsc79FJCIboLb7HT/H9qRdj6MNaZcyYz1W3WwApUybiIsUO6TqmSIaiGGy84N5q9DG3Q3
htP2WCoh5SQLdJj1w7Onk3hcK/AS2VjAAWbVvt9lwv0sEs68djMKqh1+/fchAR9RbIyjNxv8SLpa
oUpfP/SSh97UiLM6vw3G6qPJe0XzvtsePgB3QIPPW7AgoVhBM5O8y2dHNPSYi3LK2eOEQGGfiK7C
zPv9PMinkmU/PKbxFnL6qdPQT+dZg9tAZBBGWhMsYM2gHnM1/QbqKvdPz+gkx08IDUwPND80R1+V
RqrOZ266gJA2be91hHcgg5BnqEvN+nTDpcf8NK5yuprO32q4546VmC53tg5SCkkEij2oKbWFmh/W
AKP+C9rMmSP7v3FXNeaXcPJxj5JAk8Uj4HopgwT12aX3JEpNzTtom+uWWvIZPLdMAaxeQDIvHEEc
Gji2ewTd+y9t1TOxDAmxmgQ1YHFSg02vS/LYBQY6zi0qpPyYEWUfiKL5QwTp3dUg6j+2wVwAH3Cu
R8j+91frGhalvwP+V/Gcgy9l43s0fVej3FKJDFCKjyJjFjAcvzMgdo7dzr9bpb+pohcBMX1f/5Tx
M5dMwWqzebOEHqai1NvddLqi/06wxhhBZBo9go07xqBCiP2wpic/rY1Y+KGf/BEtH+uZgpRjfvmI
+P8lelO79rO9HM4CzjzrtdzP+VgZj5qKOOh4KIVJehCkYM6nR/l/V61EcO3E0Mp9Nuyk1ronHqJ1
9HjHKKzLua5raAJWyHeo2yqFPRQcsZmbzMjkfrtG00J8f94kG4G4Hqbmta2cuoF3fwtgj2EWXhIf
4lpXEoma+bmsrYcES+9Bjq3JKtk8fL0AtDeLa26QKle3W+y4gHwQoBUeOoe0fiFwtO9DbkVFvsfq
QoYZ/qv7LgsLFAugLRSXt5CuSenD2ZpjgXXkdtFmpOpVK2olUo1BizhZiad+ya/TJZ2x2M053Ki7
Fsi+LA2MD+eoTY9ueUFH1tiPsSBRktoNFHJy/HNCyZWWyxYrwfXDnuwOsfX/dcA9uSIotPrgPrke
xw2VkzNTMjdie/aXHaE1V1aO7Z/YqzSLe4INKcJt7s67RwEz52xGkvD+gHxA9YrctU7SfvYz8L2J
hAVDBNdonxA0GPDt0qipnbC58SAtjMaqQTnTSOFUZpTCsOE5/jCtaWP2Q1lN4OLI5rnHIhA/4DAf
7+G/wKGeSDM1LEeLHwLvCqXRERE4zPAKoXetKM7pRcetjt4R0unmzjzaa/WXpyvqp+krm9nVI7d/
MJr2dcw0/uCSiFPMrr/mWIRKae8jj5Lo5/6fXiqHh7jKfbOoNP6Eyl8O3hpR2Fhoc5FlsAug/49J
hSuFX2UfkaJtRWrT778M31CgIpaygxHTRkZUklSGCJKDxPVlPH0UF1QLcgVNCbttF9rSan/aqM2t
ILLJaOgeweIhzBId+2At/lh33clftcLItg/6h9djLcvRybJJKrblfbL6mZEF0SVKvK4LSzMKultV
dkCCzN+qyHgMMe5VDKSyvmnWCZT73f/H4picioq1n1GuZ8d92jMmG+/REOqypg/M6BxjfbNcC5kk
L03t9yOgiWOa89omQ7Ipj94Joj0iS7egB6PzEiWhYo+148s5R/y+T7dplaAp7aQC11pJOUILzN1Z
qr6VWrYO3Nd8/KyMGul54hoJqf7TwYVEGVxLCYC2rsvH5eQvfPB/Su79AggWdWrYzq3dx4VC9RHN
BaP0ENOB3ROCXuTQbuncmKnzL1eBUSeH7m9iBk17WX9vf0ZIgw3uCc9rUu+1IKSYRhZPslntT732
+bQGzt9KJbx5RgrcRKAuqxYjSBaYQL7EwmBU0T5UV+QGi1peqsK/qUBWnL73OkikuEHUzmrJl840
Zg9HogXvOe773gqgkd7TTEWI8qO+/OFEfSDGrbcTRmsK6qgcFhmotXlHT+NydB+nEJQDJVlwCRNA
uAvfemg59YjkwTYGC3TDrqfH3byZmzTOMnCbOMW41iSSvGFP2atXUhB/xNRCDh2+hlO36rMeDjmF
9SSlZVBNPsapPPh/StEUCGcSfv0wmHjPx3e8++pwyDxqpotxvXkitmlbgWF+BYicWa8BKcBss1x8
9+/gsSoVRb0GtTAU3QHZuBiBpHUbHsEspj1Tzro9gVIy7AK7yChw5O0rJOzNRgDmcb+4qhrF7Nyn
6AYl5/p6RKdC+z7hRm1x1k2fQZOMX1+iX6fgPSSDYJgE4ZQ2QDjVIo3iJqU+mPbz8OaYzDXsECE5
AIcwiwkOIIxN+xy+Rdj5Kg1eP3HM7ye/9gVYh7Nkqrv925HZkSU6LjNSYd10WJANqbkJt1ik62FK
aV+PAxqhoFyCwTmJWdE8pPA2JB94Tj24Sd0HlAbMcgQO/nIoeJbd8hUhu61KhHaJ09HMw+cBHATo
A/zVe+d63CwSHUYmTBsRm/B0xBAtXHnw1SUHfoLpos0MOVXU8KaN6jiLrGjOLs8laDPiOhAwOY6U
k6YNnBK9qoEmCa+lKoS6BWFVP15PQqo3mv8cnsE26WsLrq2rGxdX4NLAI6sVm9Jdo5WK0zzcikO7
nMlunvbjcOyTM4aPF32fmMKz2IJUTKLE4/b+GvfgRTcKZTeRNfEQYRV6xVww0BtAdKsntaPncjNj
O2MkYRMKlNdHBx+FGNf/x4Rj+QYASog4KhiCeODy8SAqbTTtNJLMa/R82f5JF/oujGxMRkW5UoWk
TONb2AcYuInJA6XNTNPwVmhhQsa57E8VPvkI8mXK9ELp3mNABHUQLmRg7rivJhYhDxrCoofExuUJ
WuTABRAhVabEtlFVdGq7ej61XFXy6tLW7JfpUi2/G+m6KasaRSDljXnyKCL+3GDAp0PD+D5CLLTj
G2LszEKqFhYJK4Sjkb6opfJcXVLk7uHwdPIoWe7ZWz1iFRrNm3leA4bKo+Qjq97FFAwz9NLVU186
vPnydSDwwYaLYCBb7tOOk/tHTorcmu2t2CdhipuY9dnzlyGKOOdgSImzvweHgo6+Tz27BpD/hzys
KLdxIRKF4HcA0/Vpa06aMwuf56y0KJYXqkrjQ7gcmrcL8QoH6XCUskqeq/oYMUN8Qq9gO3JfuQgR
DIDWH7lBjUAdbrqQiOGLa9FNGh19ncmmmSVL8ZvYlRd2+nQpt/ZwyYMaQTtmNH3vYnNU+Fp11+75
YLWq0408AdyDep4u0sZ2kKzwAnsdl6O6n9+rz1kyHMD43KP83qBNbg5z81BGZ9YdcvMoeZ9Hmcfk
FoAfTlRk8kZwIPp9w926czUKCO2UWyzN6G1l5lRbO/krBdysTzMxJjbk1kV/6pRk/GLyufe5pRwq
D4KbuXs91399B3kFr0h2mw3KFdWvIHktHbWTpIBU3w7UsAGszoPFO9R5PrABRQhkudqZVJEUoz5k
p8WObrO53mLenmkvs/gHarU+skPXCyW6x1fAgga6EFuc5Vzn1FX5eNh30pp4eEZ7M8hhfrhSnT2r
sgbNMkGdIxIhQ+UNErgQH1T1bIgis1qYonxG1wRWnvvSaUv+Kny3dNsLg7BVqzw5MWR/C0bZlRf3
dSSpOArWHKRLQkyNIBIQfQXh3fdsw/GcMI7yuapnpEmgtOxiwi+TntH/9jheNCx5teMbyHyGaagt
eidYJ/ugHa/jGZaX+By1WNZXZdqnwHpXa+Me+r7jrFRhgoLj9erjeSOMtTyErlOGFFPeqIndsN/r
aK0hfY/M9k+Sq5m4OrMjTJ4Pwfyo8zuCrTC3KdZ6px9FblA0xj8BC0NC9zE9Rtol+ZIIQ82PLB46
QgbKpiquS0pzoim6nb1kAUZLwzzYGaJS5EA6tdCkMukmpjQCzTSSwY0WptyA1wRfn8Mg/cjmuTki
Q6aA8jl5KSFIoosIVNPA1vi19Pv/QOUSi211KqkFeGpGpCUolUDR/gq9LfIiA0QVkEYfaf89RFBV
xg6+CKUE10oKO434ozLM9kXLiBO0H89tvAbZDZsfnApp56pndljVtfFPM78Pnu/vIFVGVHaJ1Ge/
8ex4YktOIEZzsobUfknej2wx/s+IeJJpOXpoaHFsWe21dlX4GW4yQjiMTdOEpjTaxXJnlTZNPTEF
8Gdt20+lNVBxA2WhL7WeKREeUwaFNOojfPkNaPxq/s4nXWxQiCdFqZ4kBzrrg0iwpwXWqjt9RDo6
ZFVmM6TpLw5TQyWTm9LgHYI8FSP38FF8WK8zTLZYS+yH+Xi00Yw7nJoPS9hUJ5KC5ujFOcaIE/LQ
D8OEhnSV1xdKphguatfw3mhPIRJzp/5OqmIPMaWthLMvKiXJbExek0KUjLfKEh9ik0nDpnQg/j3p
EQE6LsJt0+RTNDecP/o8JOXILjrU2T5kSZZY8/lLefrXAUE0a2ISt+ualh8+uUm0DSPPtFjEcXMD
0u42A0ZnZft6ZnGvzjHFEnkYbVi3ZPBX15f7jspY6DQPdliJblKP0I520NwKtBk4CABIEPEE7itR
g+HL8XO5C6xj4BxNwGO8b0JkjDIEsU8/mAvooENQu6xsh5Rszldmfbzqh+kCPWtFRwK3kRMjq3bZ
6kZ2Y6W8+o9Jy9f3O0R4ZDTKZy0EXPixK+Xec317IUOl1tYfKNuzd0xPFe4eSI71x8v3QgKMdBou
5yXlNGucjLpFBHUFzdLWDiT/ghweJ2niKMgWC4xTeGohnS8kbiCXRF3pnup8Xgp5+stXpoyTDxtI
rNa4qQwgogKkwF97GE10w+/oxmSoTCFiQCex4TVImx4oMEbDJ/wlcBehT0+dbRpxZzBE4EaFLQbM
KSIaEvA6YKSQ87Vdp0+43Z614is81U8Dzd+HqmDQadRz9tbcgvqJTEZNfyD/RVYk0eG/bMqV5l4s
IfO0XYMmiZYyCo5fdGYcnL5E1wMyDLbJhM2Aj+r+igMhqiICef9dR5qKjy45ZDBE10HjkfJoYzMA
AkdqD4enlVxM0+hqF7cPTGruNw3FvKV5gEy0uKZ4e2q5ojItefSfMp3mMSKns8PvFxr5gCwSuCMg
NK+jrNfWKt5xs7wWlqCkm3qULo9jPkO4H6zGABlgDO0ydePRduW08ac2AnN5sDMC7WCSa6FCJTMx
4TLMjDU6jwX19t9Jm1IQ8ABQoL3Rd2Gq2WJFVEcyjQ3nepTavKvCmi3s2YahfWA2EBSsipNltnuK
dPj/XUzlExh8Sh/u9hcb823bF/HZTaiTJViBq1+mquYIeqD1ARfuBLwjED0cMjHk5csgFYfP8uEp
rDCeaR68/atuSnjQ0Dkyzne4aEJXWq2TafkD7g6MuBPf0s32m87N31TcPJ02+YPvTRx/DQ8x42JF
XtF2ZQd63GL8S/sVXu1vE3E6bfkMgkHBqTPYzYK5OkMyXy7llZdyoUZDdaB3rZ2REdThRc3wmSzr
Jf2uw8IrisIBqHKi+JWDxjgmfgeNqByZoWa6ZBOi266rDOev6jovq2YKMbvuPm0qYYAaX8N8+uT9
OxuBD2WETaPxPbpHqsotHNnb9hiMpN8zHY20DoDpDTFeNZ7wwWpDhRhbZcEEDP6suPJPbUxhTv3S
6WoHXlPb2ky6n8aVgqNg8MR8kF3n2POafzOBwv3iS8cuUEVVFiqY50NlJZI9byfCAuPwpjfzyj1E
dZzYIOi7M7Ddhmz39+nvOkaJ2QwvQk05BE+RweRRdoEMalTGVwTsvDZXBCDDZrF/2vI/t12+KvOw
hx7EybPwJDDjLaFhZdyCrXlmeDLTCqbfROzVthYlumSbSkIUIMjqRR5VFme0GV1sGaIxi/bzjYyB
+V3mR3zdv6TRms/UkIJAUR7GAwQI5EAc429DLqMYehHAJoEOJt3Lisr0FpVKVQRDA5VLZvlQ6vKb
VBFbgZDLgW6p9DcnMWJfVRnu6oqNaVy4WQZAek3jHwGw1oLNUTR/rMP+ZbqblHm4QDxA0wyuGbZZ
SxFSC7+qrEIuoxCRr3wbXR8P6XkrEF1fOZk5jAkV7BOq8JfHVN+WmgBnCi6k+arBU9FyNJwd2TU7
9NneStccldM7xR1BnYSsj0NWP6hlALdLGjC0ygPH2E6JEw8+mHWHml+Cgfr2ZeKDt2imNcrAuR2I
ygxq3PYMOuS4qFzc7Dh06GvaXGMYb3VRB64+UPHAYGPA6DrGKy+0b+tzg/9WOLOeUp9/7+WHd2l4
+2g3ieeOg1iZtzaiFvw0p1Nz9Zmj7fxv/hk2rOa91L1lCg9MC+rjwlUzuAUyeriKTJiydpgIcAGd
h7/vzJ0M0smuwwvSutklu9L4QqW8fMKo2vKtF9VZOtDJTaZqlT0qaoSpxOk9ZjOE4v6wUSjVhRxy
lilaGZgEt6xlb9cNsGJCy7D28SjRWNzMsjuh7YmaG6/I4+6e6PMVGDkh9hSI/kVEPUhhjT0I9EeE
DVxx4S7iAQraw4H8y45Gi4xMml5q5uXxhsFavH/Jrc5eDQinj7qIoZs8urq3c18nsYkzU1c67xC0
SgOu4BiZFxFeb3rTn68O4C6KT0DEdpm5fAc/a0Do2GDXuAQZJ8jqY+1K4c66Nb1iqUgAqVNxuDmb
wE35ZNVG2ggQHlBtgkPY/Jymj5baW7/no9aIeURqcFoTppAb9WHMNIvA0nx07ajH5qu/c09QzjVE
DONR7h1UbzFitAah/Sv/xbZtatOSr8Ch86eutJsHoON/HmrUotDGtzLMQA1Xy8oqj4NFWDPLqt8y
PmYccE5Mf45qtKhaoDTl8yzVsyVQ7TBwNIBTTa7cj0/p8dKOIxJc93nQBPyN5LG1vQwABlg4TZml
B4XNIEQLpuPBRxQD+009XTWc61jryclJ4mCPiWnJ7EXFFdB0AwXRAzltnS29ZSHejBVlrj9B9Dda
wchqdnANh6HQuY+ry5/eIW87lfAlZKcP39u7f2jRf/dXXdK5pvF6UJo4Zz0YSZlcQZJQs65mtQ80
bojMEZH7zykPfOEuGty2jSZRM+MTICg59EUj7lVWq0iiul6dKaS3/IvjVxsFk+CQ4NEt2CdcF66e
edy/P2wVggY3BS88hzTUbg1ben5TQ83SyWyrGhStuQ1jMFvxdfRYvNdd6HYMB2/ldkbjVLvKHnGT
652zb9fYmF6GqoPrPwusZ1Ed00E6Tt7SaFxyoM3+lQRXOQ80LcHc+EL9BkfevjcTFLQJ8U5qD6Dv
GM/AAJ6RtdmMue9T+zEf8vZunO95fSuwNV48WoYg2/5SJJRuKE9Ap53Sb/UDY0Ng5n42ghRQJM3p
6Nh5sb/Ebr1MOuXSkvlqmsv/MhzrGVwAPGLVQIP4txlkF8HTJGFPrB0tbLURLqO7tV2ifGCssBgI
xCd3k+gWnaVIvOwAcmqyULJQnjViQjbQYC52K8PONrpyekfhMXLT4P1EfkDJfAC4muHvuyJw22gi
IkEP/R6TGEbNsxvHEf13X6J86LIrcsiBbWu4lS2bJemuV++OthhTqKLtRis/g8/tbzPlxpIE/Owt
/mpkN9zJ7X5lCkCGRpPbIgLy194pZSJj63FH+2X/LNjWTNZtWyNvngZvNk6GxYPP1R2KlZUR2fJa
2U7wXcw8LlNZSzClBvT0Pqy+1/1eLOTu8hzZK9Oc8P9D9TUN06k12MrXiiLOSs+Ii81cw+qevZkI
SHBvInQ1qAY1qgri5MJoN3u2laiIu5tvFqcYrL5Hx+QhsHaOuz3AtUoqNn/KcEp5zTNncBDkCYVV
5/a9G4Mg4JX2zny0Tnr7SIAOkv2Z6OOBaSiLSBZOCBXWbE/h4XFn0so6/ViF6cM/LkIinixSTKsk
ZFIbnuHKoAMC5C6DVxMfmy21A6fMtKD9KcE+EhXEAjsNMsltq3likLcCB4XN8XOXwis4uIdF9NlV
EYTSAeTLiPaGpAoUqJBMV4xIhCQkL1LZJ3FtUYTsLhCduqhqiZjNIT2W76sBzks7A696SkeBQAKp
QwYRDnxo4km+CVu6ERL2+V8svvw6B6MuLV0bQlN+tZGNNqbO7/ik50PZF8lnWSan1sKZdke6sj0X
7c8Lh0eYacA9KJop8MSJeSs2Oc+MV6AKBIXyysZWaQ6ULHx8eG+JrCGGnYFRoT+kKt4ByelIC4dx
C4t8rh+jHXd0abVJiv/l9JOnaprCmVgGcIG5x7YCWeqS+iHW8fiD4E7nnolEVhXLG/JMEodox111
11yoeBrpjpFvwUu5FkJSHfJe8yCrVbdyKkk3ZZtGoOythya8wxMad18qBFUS0xmUsDxV6me0R2CF
OHFXVBNUZGxx8wb5qMKjMpmHEVSUr3d9+E0qfS3mm5xTLti4mNViU02jx82np+9DnIHZ+0aX97WM
DWQHliev+37jqyYjqgnIP0ombhVAQUEhCiao9Z0YX+/wkrfEnor8Oy/aCMhVNdE9ud8Vqz0nbp5f
3qZtAypHZ7mdiEjsc7DEvkOh023bhiW7lht6DDvRxkIg0eQ4fQJ6rT7YVW9j5UbDUQNPG8c+FPok
oCzIiW+FcRqd4LofILQZ4iOBvmi/c/jELgQsPOvM4N9RiuoQVLyFl0XsiCiGio8LeemXPKd7X8Df
xz6Sx1r+1FFIgM6POhGztyFU/yR0tBcq2fWsIydYnM6C5h+UGyTU3EM1ogBYRi8OCWM7yjeyl4ZI
T7sM877kmRYHjCztIk1OI+mJzd735Yva6SwGFVE8tInOxO5EVIYZSuzxIhx7Zkzvsaa+/H4Pyl4g
18mbpovmXMZMj12LdGq7eeKKhV8auKLdh3yQJ/pGFtJ0+VyGPJejjvL8x+wq96kwgXRPm+QyNJs4
m4L4oZS2rcOQZE8JZgJofKe6VHDWMoRce4C9IbyqHNuGC9xTNgAA3487ohjvto4fAGFbYtc91bpO
Swdwm7zT8x1x88EXEafH2eYEyh0tebhmZQynDrI7h2YUJ391G0eDryZ0yC+7CaChbC7AdtIGOW9P
uFz8lXuIHtVyOx/Pru++YT70svx+LGNdwpbyEL+M1UmUGyluxVdEkoB29She8up6+wCrJNFVs9e7
rwXCJWGfbYSe5DZDrXiexg+XX8sm0/k35PAym6vX82zYrJpFwS8BtLGgAIq7KGsstLyjPdiXcMJD
cVURwDWxhZ6op1IEKJQiANPbH1K9+Neb5PLodxN9skAJLl4AMQL9mzydmUfvE4StvNFKfM4I9mn/
18uGCU+3R0Ob9iGUUwd3cWh36e1RX7qy1+iM7cczoMfUfTvq77tQFM6R0dGPh5isK0clO0bFx9a2
96PkAyxahWyLqWg+NddnYyf/1PGnqeZ8iY9uzz1Inj9uwvbut5NMltJLScE3xEzsByQ3DeTAyWWi
bzeaVdl90khuytZHeK2a/9VHKGv7qreWYjiGdPc7ZYx7LoaKTpnjnkYCwhh9PQ8PczHikGZsJqgt
GgNArDXyBWeS444wuqcznOeIwYoDhcFZGwIXVDOCAiRs5VP13uxzHvGGqqOR21ZdR2EZUrxiJF4g
5Fc9RLWjRfuGncCJsSbizg0mjHq2wvhSLAH23QnXiUCCBH5ffnDnjRqrJNSaWaKi9PTl91fTPztn
XSFhA+FLjDGgkbev5ptUdhRR6QxND5TqdAwp7pmkHTTVm6XidoWcse+1S9t9/wHTdrxNi1duGvTZ
LcDlNgCuklt3f13P+bRaysa1STcEipv6GFsgl4hmAmWO+kcLD2eQLZFnyisWwkB6+56eYYrR6qFW
G9D2MSghTQT7YZRV7Uyz48spiZBAPi3lPyZOEwa2/m5WQL/wRrQqYQBIo81uMhGabrdLizYFaNhb
7txgQEWJ4cfEjqEBwu9hhGLdl/JwfNah9y8a7fwewedrIvJuggI2kQZJ5O4u4nE+3UxtqF+wD3L1
AxSbh3KOMVaa0zMoUQjy8/7VuvgZfmoH4r9y04XvoWTVYCpJBNPGTAqpALar/+OUFOoMFsh+xjMg
/90xFXjPk9VOROUjG69Ye723ecAGp9rLRj0Qieo7Y0htJXE+EfyKlfZzqaRHcfm4oxFmRGWaIyVq
ctjJXCGZ3qQxS8cfS7ZFAM57sKRtnsgyIXYOdcBF1Z2eBWQJD6XgXWmEMJKwuoR/Lb7GKZhvMuVV
yD4rd6nMVfoDAK5p/h2yY/8mPaqw0wdEAn8ughZfMgJq+89L2I2mkDHrVs38ewf9U9Tt5/Jg/tyB
OPW5oruRCIgh6tL+nOaBmdBcsXQFyzvqtCLpjiSwWPL8tqGD5IBhbYGMiio7ZilUfZPD2ntPM8l+
12mU572jjuMbeV2yt9xcfRKbSaUjgMA5RzQRB/kWwb+K1p+Lh8L6+SBiQ/EE2wsUOWu/MNAEqHgL
dAqRDOtjkoflLWJbgj/Yj8AcRqmfrzuB2MhLkzEzZ2Dfko9YmO1SMaltv+JmHJi90zRE1rVcivGB
6pEVkR3T9GgaTeu6Z5Hrio4mr4EHOJN37Q0ok5WYJnGnKYH6PwwhmTDi0B2iXNmtlrWXpHHK8e8B
1ad1AjKvolt3jgHomLgNseYAJw9Cwv+/a0AuwglX76MzeNHGke5Pk7L/rxD0QjXtxFqcUyuNZ1sl
9SNkkitic0C+GCKUQ+Q+dipVRf3nPoW4MhnDJ850tqGfTlkFB9lsn/ZClC8gpRcxYRcoBvTC0+KA
vY7OjBjQYlchCStvxSUDOKmSp5C88iUSGVCReoy+7XowRXtkIfN99M/g8WgTIuUH+OrhrKVUEwZo
Cx/YF9owfWtMQwWL+zA0glg0KoQALrDeggLo+33Jl5m3GM9LmvPPqQL80l14NpZ1EM8ED5M0RQKw
deJBMs9p+Qb6Gnmem2rnqG1AhIDum7fGA8xIqUdsDnVPHsM89k00vOclyJjpN13AfMP38nhwOwer
gO8Ti0uQOKqNHm8uDo6wihaWd7gDW1PdpCpo68ba5xlhSRQCFzm20NS93MmYYdSKGPUBzfMQUQ+n
dF/Q0hUUA1tpNZoYJeKS/fI29Q3Gc8anFsbt4W+dc6f3Ssz0DZq04GlJ7nD/IeRNbCJxWUBITUV5
iseM/Nvfgd2oWV6ZEbEkVQxSaDhSvWpsh2HpqZkZWC3a6B/6sBkP+VNEIyF/AOvj7yCoQM0mfdgO
Ie+EiJl6U+vOiHcp/D8uQNWWnYCEiqkU4HDb9I4goOx+yheLPTAqY8Bb8wn1Y5f9HESOavoAoSbE
Z2fxPdbXzIsS/awsa413Y5uuClKNCZQmG0meykq4lVHJAI5YGLkTSyfR9oE52u75UXH8FFH3H/Og
JrTkFzyYK2EeNq0ClP91ODyYL/GiL/Ehs0TwJtX2N4eaAR3lQNY4DFhFjJpowixkSt7CRgJhuxLR
RNCpRWX4hSppHEtK6h8Tgh5iLL2sFYq4KR9PsmALCb2hhaikdvlCgT9kE1yfbLw5cNYJE4OJSvcf
a4rhlLAsUBG01LK3X5/ByKOTsREHzB3/NDUgV50XXUV/yTMiTQIPqfjImBD9eeH15NKan+w49LpL
G8mSmfV5wp6TteOyJXGsP4K2dheN9l3NUgN6USHPzx/nJSWGgOmSX985mSIAak0kOVcFst+TPEVh
ep4le1nHmMEmX7VEy00EhtEJ67IApzOqVGfxWQfIBMUHacucAWJRCsxG0Nl6ImhKKkFKksQkUPM3
KfBZBK/3RijOJE9fQsv5yOpxpqPszsuwAZaeQtrwXDA15IE7Kc0st3+zFyYDW77CCIhaFEJ2qmkK
tPeUUZsI+1iGFmJeNAPH+/yhwUg3u032tB0Yth+mL2g7s/IUJN5ry8bwQ/EthczT4ij7/Y6uZdRS
5ERkQPrYt6yJjVS+py66B1Uze3eAGkOApYVf+yXswr5fvau8alaRwVzolhFz6JcauNiXd7SaW4Ne
31q2VK+qmyRPB/Xxr2zLN2WsTIOVoelaNnd4Jfrg39LtiCeOLITYencjPEwSVkk40jUXIGCnR15S
aXBfVSxFAiPOyOuQiizzFiHYEz5Y09LayUSrC0D/7Kv+VZUBqd/7O1j3AI2J1wOYhsjHa+PpxlX/
XFPMPc8h2hie3SoP0weZHU7HSGs1AqtpA1HUiq1QITTBUgfcbrKERdcOZJ9wkAn/KKIw3dRDn+K/
Pmmmd/pfYfW7oSuSVEPLXYCbUBt/RrBAz4hYZkN2OpsfJ4+w12lKbYoYGtcj4oX0MVH9ksH/UV1q
Lf5EA2wIF2412aSsKdCSrHogpPe1+xQxGS0avp/VLpya/KnpxWbljwG9vC4S5/avMEWjltpLNZWy
nTUooRXYAo/Kj6/AQTVnkiPGvd/0hfSOmWKrpjFVoiC0cXg1YJ0s2HSHul4CJR4BrAivo9AmuraN
EhwzDZzuA3skGIYyvCFnCALy93g5dpaVyCzSCJ0BcGam7Zen4r2dY49LoKTpsgoPoMClvx97iYYc
qg0PCnQiK5zNOXddUyjHY/vaoGtee/Y5LPFeG6CJh8m6IrV+9W0RPDUkw18DWfKl34S0o30fhAYb
VUI/tg00cAGWwIcMoWQJ0Henef4aUUlznxw3Om6do3jVQYvgv5p673J2hfwFQ0RF5/0BqMiMOTdN
CNgzSESxWYTqVRRtBp6S9vA4OkeO8f/fdhnQ6ljMGFxudZsaJn0EGFNnXY93JcHwmzNylrIoL5Bt
8s+vMvUd4QbblpMU3tBjX/M9d0YfVbjU3u1pEnI+uqdWM8stbADd3rxmiRCiIXqD6UezXx01oCKu
Vt952W7tVck7jWvag5pgxfklUoTvuq+Cl8Ev6vvVLLudipJRS+Efc/e6BWzx9VRcAYAvqW9t9Won
zVQ9ru5CfED77dOgxvsix1jx9n9RIIYiaq6Y7nmoM3i8ShJ6LNxQJOans3CVCjjMs+druYkwOU0a
dpwUlTIPIv2XKyFwMP2E2tmhYT+gfPxYo9JU3QpT8v/b+fKIfqwoCiCnfh4oBB0Qo2c9qzX1Ijr2
lc3X9iwYfcX7hdBc6eLHs7EfJxsoIwtfphJ6jfOnKxXh5CHjVKsxzHjxFfwmpeQxXT/elymGAnCm
0kLmyHdhxYWiYjHMn25snKtBzVPSmfrfgmfZjeI0Bqj5o+PHtvDSHU53SvOZDQW/LHDW3oNn2iyr
LlGxfSnMmQSBNCQk5hzpqK9xMo7+itDVDlzGPaANLT8ZLSX+ELhacbsdNGq1BDTOcjdMwEeUBhvq
Llb2Z7EWy4TSOV+ne8wnftSjQ75FtQwCQUwOH48ppTTcFpM+0kV5M+94+/VYig/eXgG8I68i9U7X
GpU3gg3r1i52VKJEO3TeDocbmzoUUBsrnj2clzFgrCnRpfe+m8oan7TAxJ4yf6UpkADaEcgSi1nu
5e4b92vzg4ATMmhP/xj9KMKGkKvdlxoUYd04KCosLYlNhoV0FZu98haEveuGFgeWPD84d9HLUx0P
kavxoUmGxPQjavP8ZwdIXhpE+Bj9m9NDTI66WwsYov2JVE9nMz3S3bDUEmoqM41zJWrVZt633AGU
bNRFhrz4YIlIud4TdGLoXxGAk3kRULCOSNr7rAua5+fLh9W7PULgQm2606nksYRqj0VjFEYfVtLy
lRIn0w2HGjOgIwHWuVbhEuGkbwqibtQ5dXb4vlszMZWwnjuxWM+vkWTvZsKbKjz/eX9D7AeW/kNU
V74GyRWuUGQ72bkuIN+y+ep8uOAFZcv9aXl/lbgQWyuUJfGfrmWcPL5hyzGJ/aCCKn9n87RfJ/jv
9E9uflaewMiq5q554WYViTRQNlNhICoEgXTGUX9TcsglAFQ8d/m36sLZREuZebgSE8zzZk+pxJq6
69v5MHX6HqwSCAaMF6TWqqng987dZC3V1nPDgiGfcs6jbWR8EQoOi4o8xkOPeTkLsFinl4MAC3pH
KxHV8yvi00r8Lzi2dQPoYkm3BvmvRxcBcpSaZfzP3blyqNnygTB9QneSVunzxaAyJR3Fg4ESm5Mx
kNr7NmQ9QF4voyBDXq8V80tiH73wyrN2yoFeIG6fvPm+CoJFmmPLpAbnZM8J9JhmFHU3Wpwi6JR2
r+sA1IMzawl/HOwP7N0o4cNFQq8KlcrVxzBCtrdEFVgWCc18OiYGlYKSz0tF+yC+Ex6iknX3lUIX
nMMx9SFbuudQnXWZbGnlS7Pri9MZnb/u1wl5kP4m/qO5cqEE/+Gt1Ytnt5WJoNzVFY/rAw4/8dK7
eGITskxoaWOnR6JIxw43HWyGwF6jQ/YXB4SkNMkO1ZDxM/2yxCeUliIST3rDWybnyc5BU51mcmpR
/OaSxPTlJv5Jg79GFjtJi9BppfDJuLcc8gqm1h9P3Xydp9mnm8O5Hgk7WRCXyI2fOieAaTnVzxTh
/w4qe4+YszaY6fI7CTBaIXdRsuLqFUBLlvFHVXkl4HXaKAGvTj/Szq6qk9x3ZMHohKhA6OmGWWWv
Hp50IHmvw8yRWYaM4RzgJy5sWvdKHMhTYYVG6zvgS4PY18Pisp/scTmhbuYBL5PTbk+uNvG2NVbV
GhtEJgzyDHRTcyB2DiK041bt9MZVZ7MfU7bNaLlvtuL1mwfe8TLOAhwPfFw5+i96fcxMB1gt2pJS
3FYex1D4E5RtY0xBEgDVD58fFgkopy46OOR/G7bnQs2ri+E25cJudHFIWyClmQwewEE9UwGVQHLu
5c0IZaj9XJtPgwPt97/T021rr1PGrhXpX6/8fr7LplGukdrF1FWiQjOeIH6e/p9z2teTgQyjQtmV
dxQTR7u9AAJa/dQjQJkD6OZZpKWOlA8gtoxAUHJKhodj5RBduNC8Y81lefKlgYX1TuCukjFG4E6G
avN90ODkdGek9mioW19nky0tkr+HaqbxJdfjgf5XDOLLpmMeGRuijONPuHT9oZ1VE/penR3OCqyX
PIGRE0VPg3QL+AZlMCu/UCrGnNtazuX5dwP/MBWyA2dqSJQzJ12NfsSyTvXQ6tPZcWDadzlFD/qw
VY8It1XyyCWx647LLAalesN/RFjTOle7lrPc0t15RrO7/Xjd0Ww8/3PlBTKedWznd31in0Y15GJX
+aioqFdj5Whp6lXBFSYM2Phd00ibzjhisTWWKrCIb3OjU5KaF+Xb5KUpk9YMx7PnzDs3WKY+4YaR
238sWgEbKnQMlQ6i+bk51tLB2wXtLOdKUdWZ2LxoTGKGAD2rkR/JHTkkz/0oPfSjTTgVfah+bv9J
GUGB9aNFbIiwVn854WoxMtUDriq53/VsG6zAMOVHecv7KgwiKXUaTwPdiKrzXQWMjpUxPh2db+/U
YtrTOxLD3qHIoiUgvMwjmlRvfLEhbhib6ymSuatoxNTdTFkcPGv0AvO/En6oVDJkIfJkOnPxJLO9
Yb+3JHYR2ls44oyLP1+2NmaWSD1war4SNcmpViYegdkINWKGpGEDGGkg1OwKuHj1ITyInv9NTE4W
2O9LzuQItp+l5qqrQHBFXWyJNbiL9AAWFWCod4Uqm7RFSOhWj0xAiMeR318bcB1YflZxjYLIaCLT
pyUSgE8+0BLyupQX9WNMNjlXlYi6eGYKI46gfQbxHeJFX4amuBkYgUkQPJ9A/n9S0urh5HX/SvlM
o1KLT8xLSxjNMnk4XcjDq6L6Dms44vA3c7p38QwkUSiHv2IevrgL+nK9utd1vPRncHah6S3A+ig4
2gw1a4+2e2FMTfo19DsRvbrCiVM8EaDaE7MwzMT4yFrTW5v35+6VZPOcNCBJdUOY5Y9f5Hcsy3Sj
vEAc81ITdHciP1z4q/hN9mBIhAf7u0mRt0GUDE7PMqjz0sJGQOZhaLMLlLR6Zdexq+AXm7xPGWWQ
/H9GTI5kvNIYjubWRGthRzCoumQ1xb4EaienRimEIUNcelOhj+qqRoALIrVPrkDW757+3w56t8t4
S5dSsj/99LEQUJ/REzApLubZxZSurePDmvEzSwri5WXyCqzwWqKRNlC7oLTtWM5lksiPdLNta6UZ
NYaHPfaP2Y4FIfbigJPAaJb3DPyuR6aGXuK/K4iRe6g6U4royvITl1Y4lc5d/Q08AAtru+irDpXE
3KXVZrNEqaVQX+IEXwvkdi6t8/BBBk9uqIdF2gGswuOt/oHw1U2SwDGTOS0QD7qcvUtMl7Ulrde2
hIh9Gdiedwb3+HWdyx15pt1iGclRqFsqP8bBIHj3k1foq7aXRcqH2hKZSl24gBgpnDQlqBtZIFmE
T10oEEgUVIGVC4Y0gKn1y8FHPwNf/C7m6pXxAEll2einXuOUtl1JvBSIZM94Y+FTu7nk9wm4cEB0
OXFY6PkbEwUHh8FHsAfCNc7/zkQxgbsqUeHa9Aj0h5JKav+8s1/lOcLJ5/12W1KsxTLXOymE2yYZ
ugttdy8XJ6j4lNFEbnPd32b8XDnqY1h0nugIP95gOx1zSSVBMLw+tIZ5i1YCceOmyyffFPYgpHCO
ym1Gtgr6+ftRjPfQptI+xFcgGCbWZ1Px99hdXVMr3BJiNTuvyRoAsEL+AUVAromFzaNSEon5lIQ6
1LrGPat0ycU7O7fcLn8P/7zF8o1iStk3aks4hduwL28oTJ2Dar42qVWlMO5R7cERvGfKCK79hIB8
KtsMcFaxatqwYXX/j2CuNkCNvPVdCG/GDZVung2nlOvqIZ+wbtDZ5HK6u3S98Ar5ZhH9Hw8fU2O+
Z845BmY8FL9W2uNJcZ+WtkJosNTTc4qVf/Jl3FkSMdCnTlf1ZZi/ffqVv6N+qztrF1TOB4rq3/MX
H3RfeI9Jx84qiLTSNKXAdUFGKfBp6fbuHssJiTDVDtgiWjVPRNOX+yTsAyaq1RwCRJIps4i5IBrg
NsmbXJsQRrWm51a0BfF2jqIsy95+FhCLnxYJIHamIu2Y9cjPaLiDFpcc2WD6QzJ2vPhQRIp9hlTw
5XwqeyNWCtEJGFA5P4Wq0kQu4ie9NhPGHATbhPMmQaTM2i/1ycj+HVDIdq0EnPZ1FZXeQJ9tNamx
yVzX1IdRR10yjfEHy2/9ytjOX9UCBeHiwhdB+tf+FmDVY2ihTVCXD+tb7YwH2NZo9zpLR+4a3OCQ
sGfCa6zExOWLYGCH+qfFuOE3cldEoO5xKANH0rN6gBvk2DWoI01/lxQClwyO3bUBtGPrIpVgeTjR
Hq592GmiBtqB5TeXrWL6H23gN9X4th3HMaXhr/BwGN9jFHDfHz3bM4mSRs7J8UjRuLhSVKWSRLw8
QdU1DVe/GkVvQDxy/UA6Sog9JLOtljhVr6qjAhpwSHeAL+UV292ZdoobaSVL9sNxzKo7F6NBfNPp
BWkqHBRP1Q2pJDJjqu8dNumtc1/QEB/vXAWPopwwwVv+NLUYTm+8qkJElym6UcfrOSx2LmOTLBnb
3Mc3tPWDoujzepmpTyP13IJoQ7JqhZnZ1CCkbmwFOV641J3PqDdvCaStK229T//YLRwPR00PxF+s
0M4wl66tJYlQKJ9s61paLaf8nIqCcbAuJVeGW6IiTq5QN6dbOhRtiiSEOZdvs3eSJkAq3I8ts0kw
mxS9M0Rzrnbw6uJSJ3kbfooseSd8vkJwPOujFR68sgnjBW44+0abHuTTP+KgzUVwOHouCNJ62LVS
YuEVDnXZJZ/v1RqhSPSorxEJ+UqwMup6J2VNGgqTck/CYUQlV8cR4KbGtqtzAQLMO6uF0ClIBbCb
b6cyiTaF7NwN0UzS1xpKwzKzNdC8bvFjcF6IAi6J3CeXHhDn8x0o9VR4sz0ak23BuBxSQrnyKJAB
qsxw3foNWRPE2c6YOdPWKlvQWieW7pg/reLVfGYVWoOI7QEb+uHibvvvcej1kT7IammrfCmW4DGJ
FbZPvTokdbl4SWDTErXo8o9/mSqOg20RmlXsMHLbldEJOp0pKs3UjqoCz8O9qN+aFVEfk7anj7q/
SoaijYVhh1Ukjs1m8G0JEdvIBubQij6e4iDsrOntPwyiFDBHXaQUNcoS2ScQ70DDfiBDoj2dk3Vc
2mkrLGh7EpiVdBh8XspqfgXZS5u1kCwly7gfd1yyyXwwkHobw8lCVk+qwBqJUIB0c0dNtT9qh120
XlsizQbZUdcK/BRhEYIU3HWnJGiZt7HRYYRFm1pnZ11bkA01RbmZQwgpKvDmZoo9NNrXOdpP+ziR
1Pcz9SqEdlybig0XC9bnHMxrp6+2T3bGZ9YuNtTq3/WiD46EXoknmlsN9fSJNCrZyg8qioQM3+mi
HdFKuyS3gCUe1sOonQuEuJCMg8X5eFU+0/o6EdxjYrOJy8tsvintHY/NL2sdbtASvBW3XzjJEvt4
gGPVlar7ka84XkjyHWnT9QrYH2DgosPbKjlHnFs9ru2JkBWa+ivRyNOEfO3yzFBSNI5HEGqs+WeD
9oebpGzWVMwudK1wj83JcG5ndHuNaZv+LHOu5fj3MvEGIeZMAxKYQZzYWrE1Rl8kIpnrfzd+H0Bw
P2bn1W/r0RQw2cszgjngYEmZlLo5/LFefOi/K/2wTxtzjCPtPdMiUBVzWX0UPshVCKWhfnGY9c+t
YtPeB6wpWdrC1auyX3TUnjuCPRg3pfEvqElEYFseRdoLqJlgygkAUBuhO6+Wf4N3c+h3sSwqVxnt
3ZyTS9HYLTDWfJnhvCfYKb78D5gzQhtGIEKUPsTP9QIS8TgnoOVCWIEZduwmz9xJVtEzXAdv/WYA
PSxnLCUUXL2vptcxhYbvXbjBJx7Q18bVCA2iSkLvQnRBmRMjOqNv0iN+okCx5Cfypt4FXrIErErq
MmIktRul9G14MCc8fOJUPo6Rjln2twEAHc2s6NoEjw5sc3IgMgTwoOjR80mzV1w77lVLRjyZXZvn
UfcSt8OZd9tFHw02CmJc99Pi03NYb6mNDC3QQl2OWEj5UGQ6Q8ADW1U2LshqEYXyDztvL7oAJJ4h
nGfvpNyPL++jnxjhot8aalatfb+GrhzMP7B8aIr+SDSZbBdwM4TSzdJepaaBxVgDxytAfVDgDlYU
w/uyyfkVrcnKhuMuwHHNx8wf5jiTqhU34stFHmhHo5pjipFADi1NEY6ZZCeq9Y4FbG/llJEJfEvB
WhRk1s/CHIH+/eggyWi2edZvDpcoUY8AdcA0gz/ZdK7RxRH3sWE6QMfaHpjCW7rwHwu3C1Gur6Kl
qXbqVf103xRfKOO9lIKXkYBf5nAWjdXt1taklRRFKz+2qHKoZRsGuvWLtq7qcxLxId5ln6xizWfy
s2sK9uNmIwK8fYuQanj1QgUqaeuKZ/4ugVyyE8zUj1lTAyUgFCk5oAIA5sdchMtSCwOnViiPYJQ0
iNfaj7gUrvMPHSx37CzJIquja+YpAexKf8pDrKkyGyBxh4P/S/ToKENokk2/P+c9RguTeZ9JoO5v
nyKXwMv+G0p2yHU9h1UbcyQZs23oE4dxo61QlCp6eWwcHUaUu2j1mIqFMNtRCJkgMneoC2p/6l9C
5qeN8x8zmBrceqUGoI3upS1jjtDJDBP7tWFGvMk75zBC3fmdIP2Qi3gmRGvuRjssga5zLCjWO0eA
XqoynjLLO8hewkfzZdEIoGGkNRPzEIiDhR3QCYIIA+b8hs1+aDbITvhJEAiUu+K9vMksdk9iIRkt
diLo8M15hXl4//VU1GXi+9hmCVRGsThll44+eVjhWj7Oy58qi0logQcTM2GeKMy7XyGshuGps/ov
+0nBUUC70IbIGrPVylBVxuAPjDcZ7/zhh0b5LH3voohtsXtFTyh01flh35CTCGotpM51wXicJIoz
m4kLfmp/9lj63hCsKWz8H5rWtNAx/m2emxm4BP/ZOTDagYf18Zy0DMKV7pLimBtxLhKsI1+fgmIo
2mXlefGPlcTIPb/sqiPwG7dKqzX7uwl1sa0f0O084kM9HnDIC5i86/83e7ZwspElnhRqfAtzfC4H
885Fb/nEsGW6FFFFNt1kuWrVNdkrI/l7COUbOUaDVlln2LktIAd3Qi6oW2O+yG+d1usJ+YyPojId
aOPfVqXNoZwdle2oE8LvWY0rn+P4lBVRwCgfM6wguv6UfEekmUtN49t8qegzxOBsxSQQHWMvLJNq
lPTXeChRyI9J0Jz3ANIREI/+q73vonb4RsNouuUM3eE/c9Omi8Ktovwmq7qBa/OH6/YxbH+/F8JU
ZH9wNzQkXkzVeM4wTQW5HCpO1FN+lA6/YqHTUXEjhaQxoMMIuFYdRM/1GEWl2AeYtKKhhuZ5pabw
2yn9SNpOnqpGq22zNkjJ4RDOZPI2sntYJml1lShGw0bUkLYRWMTbyI2LTQyPFg0vjRT0YTWkapm2
vUNd1a0WcwCzXkIuqEo7y7TeFDu/CXX3eS1TNRlEAmjlpZlNbEmnO9Sqw1cVYA9J7T7g64T5ML1P
7Ufj3RWrFbNbqLYfVDpBe1IbWgv1lhqu4F0aTEcqGzo4HAsueqJixYQRt7gqVfCbY7Q5tDh5JZk4
H8aW03yxm3MuKMlcJFkgG6oPn4BYFljWzxZkZp8YzuRAyrWBKpdtkYZePEteETyH1gWv3u4RZo9U
6eZYEP95K4E2e+PdPAz+J+169s3FTPO+JCmRR1WoR4QTs14w57vmfLnZnSIp8iBtK5oG/p7WrIoO
OWPoI5b/XJQWKn0abgyZ5gpLlGTA+CN+ag5nhxdYcg6H6UQAHJqhd6NvCgl/3XANttOnWiuBvytb
Ria3jtiJTGTha5JcVhGfo0iU4BbuJ4onoH2C0GtZMc8vNYldkdp/2BwaZ4pL4MYXCOD4F783/kzo
x3taPHQmF1OuC7rT0qV1zbkmrmJPTwkyxKo6kazaqLUfeDTuo9uLfQS9PXlKLpAvZ18if742GhGd
GbU8Ml5D9VtKxbgca57wAgPFzrkRkFG9Yjp4jiz16Ro1agtO6h4hJ+BjX7yn8DE6HcQAMXd9NFIg
n/iGgrWK0f3uv7j1DjRztIfZgrAKDGTzTGNSPuo/pwJSgYA7TAKj6O5gaAkdcRfINWw9tgdULQg/
xTkyKBvBErMeeRZiu1X9UfdppOfK1Y0Bqp105waUVSD+2KKN8Pr644ygGtYPL2VocS56F3kyHJ04
yx6oKUK/Vq0xnd2o+DW5vADhRFOBxxn9JvHzeTHPoHXYycZjIKciMSAxdXnnQm2WNFbW1Sy4Y17Q
bmPL4bKarfHDBi4OuXhjhIHk/beYxk/7rVPY4cjDSsVDx+XEiRy/gRrUysP/vmp7pJ+Vc3HGd55T
ILYy2sxLAK4cO+Mj6hw1vrxtHlJrTq1zVR1aM6ocjml5V5dh4oadAzTmS4jqUZNGZNp07VQjzZDs
5EWVNZ443ohCjJRCRXb+6cG5BHrA9I5W4syrIfh24tRKMovy2dlbzQufHRBD+iAFZEEGaxLfP0eI
BgzSPEVBto96A4JymIcEpI9Sr9fBeT395mJerbcgqTpVE5m2BIvzi6HVWKWPK5kQExDdktKf7njd
GQHiyatv7cl58dAuhvUYilG25FWW3BgYMTuNpGbVn46Zl7LyW6rrk+c9mHSIhiL3d+zMJ8pySAiq
f+/Ik4fbn85O8xox3MbsKim+/+SWFoyQ5Z/6f3fFJg8mfT80+newfOPA7UwUJa8aySGB9tFfqIc4
booELSi1ogEMHsmGGIduYyZ2WhNO8y4csf0zENV/q1p2R6kXF2WpwLMRkqL7is8uRvsFzTQ66zPD
eRo7kIQqTXNfgwAqfG7A01ePzsgOkegnOdQF1nEKUjn9NzCU53longubtrlPmzVkrwQoAXTVUupE
6B+tZrn/cfUEvgzJB/UjhGkYPZ+LkyUQ8Ehx8vkQbXT6KWGk9u7kmxcSJNub2ZnehAmLQgnX9q3c
VoFJ4qx4+EmcyClc4fusi4/5T+zIISgsv6srOHtkpI1jhiN8/fJpobETJl/sczJoxQAL4ZJVWJcv
vcItc9SKLgpYkvrBo79ezKbW+prJGglbXxLK44DgyklS4Cr53aSN2Arvxme+IuXtp5An4a/++FK9
mKSDidBGJwHrDESRVdpF3jbzU3noFSTbYsRyHd/T6EVoFLwiFCTAkubGbNMT2aGpDYmRH9KBVdbc
TXKIZMrCAxNKbxMYM+ts8vpeaR0wX6tlsWe8wA/rB8lmE9Ga7kd0DTh17NETNN3jzDAsqK27rFTZ
yq3oU1EqqwLsTH1zhJdvmjagRi2/oZ/KY9Z+XMgEHelmGcSTkAtCe6x86pD6VyPOcQtG40XP9ioz
GldYMvNkO1VGc09jzbqxLLVaG78PBLAopr0/YfkHEDCkPoPShfeNm8a/WaEV6OJvpGR7MDTEn/CZ
m61GuH9CxhBqt2HvxTySPGQWBB5SwreytCfORfWNjsUcvmCV+hZ8CFt4PqZk7hOoyCltNnRWrz37
uvU9QUv18oOmqwIb6HJT1KTEJqsY+dDcitLvBEzUA4TfmVOkgHWQkEb2rO5BYfd4yUzmJuCVq54p
DBxm+gsVfO4vHzG1guheAQhYwWHFwL8EZGDB5N0xhQUIRvOrf5GYfqrsEE385WA/zhfgP8bjPQ2K
Y/uzB7Q06uU6K8M328QLML7HYV/pJK7zd+keQnkOUTrOXzmUDuwgE+ab+SZEV7esAEQwZBDe5Z0N
CoRpPyHiDLLsEknc2yKaYxOkq5/nD5dtTu/uC88f5TmE/8T1amjzlAsnePtoq8nhtsJupVf8O2DI
meSveDKhDr5B4dSK0Wzs16xYhpoWmgvTkTYiZdbYHUb+BjdqUR4ZE4NlL65jTG6//m9jrCbN0OwF
A4I1GC1gXQr5nBuLaJcujVOLAXmBscco0Qti5perqqg9dx/f2ESjy9cYfmJnfh4Vzr9RnrspsnpT
xxojC4J2GaDX4QcWkxRQTAtQZAmS/lagg/1OYWqExBwZu6FYHBHz7D8+nQcgVcQnDXsOHjirglyH
ZqvV5pGD9EC6dplsWUqYMcjOoSW4FzNal+lSy1CklkaNFEnkgjLPs+8h4n7iN/iT2emIUXcHhetY
nYtZHkzk/vr1lX0RE0NPx6DzdV55oo4VaCXLm+TNSAnZekl3kWQnJBALtB+JpUt+mYug2OeqrCKC
dNyYQmZL7VmiB4UqR9QBw9yJct+gA/Skw+AX/f8Z7CVifCsLwgSuqifkczWVnDARzTQqVtMzcPVS
1vGsVeTaRf+hJz1wX7P1eqkDCuAYdhqXogl7+C+iAdsYyIbGSGVPCyWw3pjIbYZ/mAYhn5Pd89y/
AMxfdjzcggAX/M+DTNCy8HzDp0IhhE29Qa/TVN/iD+vn00Id5L4WxaVlKZHgJrU2T06P6G1x6zyH
F+6ARLqoOmfwYnD+p8NYmQxmfjcbYEI8+CpJrsdytgZ6liw/fXHmLaZshJjxAXucFAvRmdKdMVSU
17IZl9lkHCcrz+wXZAAAJYNFNN9geDMpMiWIqY4/AoQ1pdSEThSJI26rzXc8Wd2uLfzaQg1UfFy6
dYD22kPpdS8oMivHdMxjJuW9NaXqkM9gBbl7fxKgDnNHYOmOcsYAxDco3xG9NPGDYAS+q9WjZ2P6
qRp1mdH9dsJLZUWxPzTZqXhaazqQC7kZzKwo9tVct+uitX1YSIWDtpWFqoBxNNEZnSzjlXWDapPs
GgpSUe+FjsSf7CtgAz98GmLjUKgS+/GUK4R4kWeyKi0GGOiq/fjlkZ1Q2r5EeGWX/WGtnpFKGBiP
UmYvOpZG177GHwWs1E3+Q5sasYTbTqu2KSWh8hrSr6B7+M2GPdDZe+7BbvklIpWy4TTkkZZLANjM
DxlKLGpUBWUeTRAiQ3Rd7fR6e/froL6jKh34HcyiJ0n/UHeCA4spYqpAIFLvoyvGDZfgM3h9ep82
MPKWuQk7MjLlaik8bFD1ZAKKW1EhcVmUlmlhsWkkjXiUedUNgAHdgYNZo5/Tn4FGJvJi2/WglFiL
avcsvSKSR1nufTT6Uudmnaa46xQy9cmwKPrFOwS3NDuQF3Z7RWgb0SpStwT5NQ9uxW+3uw1MIQid
HtM01zI2AvPCZdBDMH5xqRfFDPwR9tLs/ITu8Zk/1FJ6mI3RbzQ4vZ0tTSG2DmJGlajoTfm0kRWP
gi5FdDBE95aEyXFGkOcrrPSFo1UEPXGcy3QbBTo9XbcGivTkuk8N+wKM9efm9SJBlXL+2KIQ7978
EhxBc5bCNrO9tm6Yct9OZRGq5tjHmczVJAglutmvqRm4Pdkrdon1Ioe21hg9btpG48LCHiYR3Dxu
NWT/Xj8ya+Eyui5ck6XtISOONReGwed/sdpDVsLiaUoTH26slvVoOkWMa2WeupJV5QhcILBdKcXR
Errnf/jhkinKrzhFUHrT2D35Ja5yMQAXO8yUc7FuI8Sld05mCHzMwHowWyrnmHgSBpET4GRBDvXc
qYa8wxhEW+MOhkqneS4cwF528PgaapC9/QdfoQWUxhBLRn0SU7EuxlcibwvLON+tBuN39K/I0XG/
/UaYIMBBdINM19kDcmzWJOG3rQYuej5ip7Sre/enpKLpFSfMPGNELfvfMElj4RJknBgytV7ja8MF
fqHww25XPP+XjyBarNMegM8ed2Xa9ws13fbM0fKQJ69BwMJAIMSgPwisSHlaQ0w7Y+oc1aiL+qXk
04HuPsuMFEjTkKIy4L+wOSHJHac0yBKdrATjUOPx/ZMZoqXhMLzf0+L7VwebluuRgOFFKeF3MW+C
XEHX2YkiI576EpDM/ODGAMBgrG7JgHJzl44rKHF7Bgo48MlgGMvtyts/ogWV17VI+p7ByyKXBbQw
acuD+M+WHrVOvcNuoQDx/EYGDgsYhnBf7wl1rCJMlLewTaq2R2hPnwTkPQKdNQIHADQqTfKGJdsG
zwcX0SRkIGFRX/sPseMrqOPj/YzTEYUdqi98lXwyMp3+XlF+0EZ0C4LsexFtc7BjW0EdWDJw82Vu
0PklmOnkDZxAAd5hmmOhy6FvwGXpq/WHbNLNDG2f8mD0fY0a7Yk4jccm/2js89NUxW610eHX+Afe
HmWQxdT+grKdLejf66z8qbcIrPyoY+TUha7OKYGgPYOatMj+I78uGUShtZOgRI+txiBjVV2AobUm
Ux6G5qCPpSd7XK2ZeD1Nm8U8ymDNdiQti2uc+hK2L7K58syUMAcL5heQ0zaDHDacgUz0iKFNXi5t
isy0v6zAqmOPhbd7GOlxugIYQ9rZIcwFKEkBKUDw0MkwKm0B0d3OM4rYAlZb9YfMcEbDKjLyJKZu
KTg7idUSBtIO4IJK/TgJRHL3ghOSGTr6RNbQ55BPqdrWCYv995Xk5WR5A+Wk6HsXtg+vfZlSGcRT
86Kf2DGrXQQlaJi128pIhaNlOnGVjzTVd9FCoy5quJJbitmvTWc93GbYMIRpn/ZV3Cbmzoi45KGc
JePRnW0ymkKE4GwJ090liviGYUmCjmgIL6A72PYAqOWuBeHeYXy4jFQ8RZYUXIvjY+/c56iVEh41
+rgYsiMGDHS1niaawv3ZjJV7f7O28Mife9cplizpVFOuASLrNhdK9VGBp8LEspXNXAHStagNDHTi
9H8JEkSnTQpAkK9exvHx+4al3NzlS5i47IQbhEUoNyL6HNw+pQlsCn1kSShCo5Mub0SbV0tSMuhG
PE1pZOlQdBP2DIRKdHEXC9AWn9IQD0twFBlCUnvQ8lBQdkVp+ufE7Q7kXNMiLhNL8Zk1CbE4ZZyN
2QOOhVREY1R5mVlqdNyisBHnwrFCIb+VldHkPEW2+JEo/blwa9pKx7g8jvxO6FaKAe0b2cJF7rZh
WKaMzn7ATpFYyaG2P+s33SzUL4mdXHSAmiYcXKjzjbigQGtqJnGs2WvX0oeXh1Is2Kl3Fnd1rW9f
BPfJ+IM0LnSJ832rR8VeifORNFhHGMoa97mQ8A+bmbg8Vq9yU4Iqm72L0B5TWSop7GcHo9S2on9y
e1MRyPaT8vLyIRc2WCNR/vA+QzftuklOGH4kJOOhz6X1jVuDI+ryIHzJmMINdbzCd4CZcX8zIise
nBre2efXarRMjjAeBk2i6c5p/ce3zogVjHd+ZJrvjsgiVcOFQGa9RNZ6mhQa5vUOl4bkSd9/zoNw
5cjTGUbDMuagLw5Pa22qamfrTjWtF0/qNNdVLCxJ1VjDsqKWfxrvI7l7n1E672mR+x3eGmPzBuBC
UeimHuVpQVOxcHpwUVw7OLLdSXiw28m/Jy6btSdYSYK3y3LB7zBt9xLwibV1Lb6X3pTPOaxYtynp
Ig49Rm+YNFabDhQVbtmhK2sGBePYkYT918f6SrHB6x8SWAxePjeGTOCyJbszr37a5dd4d5Vskgy5
yedjEXnXoAK12a6k6Ui0ratVPZvfMzLqYqqV9xTCqysNqMwVF+5HogxWNshHFW3kpfq+QDd63WKr
hXXnWBf65mk7pp6Ey2Hzs1fXRgOWcaz/kQxVX2TViZeJa0ZIs372SL6nkyOjOOwU+aGm4sADbduP
KwK+3hWDCO1Bsmk7GJslyID3O3I1XmmoWt6e8Ku5y16tT8pFsIqTol95+2QwHPeouYhisQw7SOrE
KiUvZ8sspdUV2Cvqc1Ov07ROABPzuWEWMxc2ZIx8gYYgLfvPIyQgT/n3Eyp0Nxc4nV9X+mXG+j/9
Q8zCshZQ+68WgwKInNjl4ZsmbHEhUTAI8R+tQQynUriha/P0wxHnBzohkByxqhhTQbQhvN+bnKOs
MCTeo9hxPKXsL/RQBvkUh0FoNglX42qQyNhuge1ZAEuhz8AmYSIM6g9S+Q694g6Xh4cBO/p/m1fz
FoksFlSZ/L6Djw+UIfGa1APWTyxi5/dBM5S9Unrc+xclg+E099ApLbWtIK+i/6O1OHx+Tm0/q+xv
HvSVGebhOjdbVO6yIeqjw2G4uQFwkuRQ+HL4FIgxbJ/bNZ0BGZ2E1Rt9l5y1rAJSC2wbHPkc7iem
4660jBb12cFkivxCafTQjqsay3x6Lpbv2+N8loJWspdCWKd7I54rVza9pNUyb3FzO+46QuhbFY/s
e5xVV2CVl0w2J1S2lvk+G2DzuokC76m8Iy2Wk/FYjpPbpUeJ7kin/ZFDaE2G3Y9IH8OFxqz53Q8K
B9aE3i16n/B1SCevvlUv8IOHqMFCK+S/BJ0QCRG87t62KsFSKLBq6Eim6B9+Qb/4tfOfcxOLQY/y
Moe5DQM43LHl6pCJzT5aIjVSwUm+1Z7jibEoirRZrvkHYtVYf/+VUg1nTwjxh8XTMzU4e1Viag8O
i953xSmUKQWnp0VZ06ePeO/79Db4komajH0TNIydyiY6SqQC3I/VNrcYphsOgQKkiqyD3oGveZmV
eLrcSv+jd7+efxSZnvOWiIGsSXc52FO90eD4jmfOF4wKnzc/aXA7gAoyn4OYh1IgxYYpZeJv7Ose
fwcrjMb8VY5bC8ZeREVTl1rcLg+kjOdQPTbrkrpdDlGh8Tu3+9h9uqo246fYsPizO8wEhn9qR8++
gB/yb58GLmvyjNv7z0oO9fFN7jWyTvlGCfiHAHVzRnxjCMRxNzkCs+87rvKpObrra9zgqYoV51cq
Ynr35GEkaVy/wlP4G2BlLV7NvWDIQM10zncysnHdoJUGhxPG0izJVtxiFTn4wRt8TQeFXqR4GsCC
xIM9GybUp2XlSKDr2Az52JwQtEZ33rpMKD/BaAWffNUeOVci9dWK3PAJpL/+7kWLAhPlaUqO7db7
FwlypJ2mxw0qNSq4YAIf9A5UuSGGn79olLeym1Pl8prIZcFwba1ULIsBhH3KY2D81gEhFYjCaKy7
8FPcC/VLjczCjG79zIwZ4GOga1PBeNBmMXEEyx42jSvLMAnp9WmqvTqgjGHSCk7tZI7CLGtv62X3
0MJczQ/x7Yr4Hoss6D0tDwv6t9/3k6TtAi9MSqGzua0swNqyV2rBf6zuwa98H1//TdPnhIKwWZUr
ZRCWiljunK3jBioOybZtGLzDRoKOs9SV9/H36zknTmLznuoD1Km5SE6e7pd32BBB68VvLDPxWZnl
ceYHcouYijz7n64RdzQTott6Uf40v3FHpmYBU2vxAbYlCDNcNBP6LNQzymx3mBSCH9GPpj3dx+xh
DpJWYvTVH4N0vTNCsuE7bSQxQN5ytzXdbFTlHZcBUkNqKOouDBfMHaVFNH3F/zYdy7l03PaISGkj
CrVgcRhSIEbemeaELndQriRkBg2aeN2dML8/fDpo4NSBYqZp6tRnNFdTfzU0OmM7rv9tietjZs9I
9dY2cdqujccJJKLO9+Aq4zTwr1nX/3cEodAtUnszdjbm/x9A23M/8xzNrHixPzIey0RbuaUP9WVB
LJmieYbjxvYY3zvJR7vdSnBXmXel5MetLNivI3z0DT7Tc7dahf8O7w+VaVRW46v91dc+VIKSQJVG
R+ZVRtGG0oeUPsCxNRQxOE9BAnyD0kZC9BQXVVAfYjE83AG8iT3ywRQWa036l5Okyn6AnrW7elj9
ALhnXYs0ZkplKSuMuGrxrok+dfxKpFPDPyasMOo21AbQ+ozFWa/dtr/g+nYs9iWa1jrKxn2W8hxz
QuSN+K51gNaWjBkruRRtyR2aVO5b7lbE38M7vj7TF81+/XsLAUiTzi3+YJbTBaU3tOG//+jiQUoB
n3OjxGacuL++qS3sQXEjd6HrKnIKZYqu07jJsKWPpcYF389vOpgkEdWJ6oBhFTBAr5yu9Tw4LvMA
7ktGhcOEFlWQ/qV2U2XhGQY616R+wyAGdmLnBHjcHSuTLwAzdUDhGzp8EoRvswWHY7MaID4GK/24
RLY3hsO07/E+aVALuDu58fZvyr/cpa36vgUV5bVQE7CFbbv520ClyBeGUNbOC+W7ETieRGIll034
pZSPCoarDNaKiAODO0pjAYsWozjb4lYxuU3e0iyt50BOo3QFxrpVTOIQTNNNXksM/xCkG5OANrX+
GWg3eFncI9hJb3Hz5VTBucJOzAOTedLK9bwLQMVp6MeJ4CaD5tGsWEyD32Vwh0oTzg1PRHht1CRW
fbIN3OFUUTs/HLbidiigASYPI2ZRGlp/umUR/RR6X43DtrkbV34EmcMczBo8EK8OmqwFKwJYGwii
x+pgiGJ3a74hHIIqqYzLYTLL3XxMnCjtd6MOAdQQmF8gVN6tO3vux5e7uYXgcTSIbay1/iHnleMm
YVtTHJ3KTQshdx+CcTJjt4h3t+U94vZ5MUGOSfExBEja+CqqslFe0YBdWGdfrBOtkwrbNFYTpuEY
hyPzClnHP678VGlMgNqgSScwfewfLJSB+eOOF0TUi3fIQcgmXqUOVOD3+sHePSwiCT39AYvMljar
rbJIj8ruANNpZ7apbx78CjhbtbvZxBqWVlR7zPRPj8+5WSGlufxxUGtA2WT11PSJzuTiVcT6xLkD
bQxus6K8HKBQv4k12JA8TeE2HnPP0CTpZfFKGtgWy+Ryu1Np9iLNzzvbo8dEpAwmGKJ/eUN7game
4Gql1w0nGls1csVuLSqPjYbQaOleE+CjOXxFywqZqHcmq9k3rqUlRXqtoD78Cx4tygZ9f0/KZGwp
IWrXU5nkhaE6/qnSCcTUoLRKdd812H1fozuRB2MLPqWXHu7X1mq9RP+vQplB2ukC0DSJbH6/nS0j
QIVNgamwUtT+LQbGU0GvQCRG06ejIIjNoqNWU454Oa5KIwTBN4NbPpq2Z+Aasos7fkFA6+fuMtk2
T1yJLYkOXH3IGiyDwlmrPndY7I4S2a/snWZVKRd/TyA25KPnLdRGgvxgRpOZ7bfLcs644VZq4t+x
tWlY9UVNfke7/Vcve8bfKsQfJOkyTWyRbZXnqbtfCtw4+ScGX5gZKU0HC3J0Ho47mkYFoNu5EKDw
31kq2lbamv3e3tOAH6jkOUQxtfKzxyv8J7Lwb1ntz6WeehT06Y70OU36FmwUadtq8DXBW9qDOLtN
2kDjdK75PGL17lav9V1xcR77SgeW6khLofMNEKLoja5NX35xIx50UO6tZOOurw5NX8SEaTYFxjlE
zLiHEXatDBnthEcF7Egt+8QKw/EsDo0/rohc9nUxoAN0Zpj/bc3trbkktOK8yjBE4saCNg7fwnR7
Sg3ow56G3XmWxprwDe60wT/ybqjHqVGKxmq+PZHKOnOsuD7dd+1TsXyBl5NIzqhioz6C4WtVN1NX
xzP+XNkWoZJJRADoYrds3dMeUIcaduFG4aNHd74ThZDaxSR/b6LrWu/tOZGFj3le87/CXXCq1uaE
JQXIBuQWGceVXeLpcM++Gd4Cy7ZyKB1q1HMsx/uiqDOLwoFKMtMSA0fTBaxkyyTYc9qdkIFl7dp7
K6byv6sU4gQ4mMbpnqKRp2J9OfbdOvhZw1Ny63EEXBxAj/MxrS9vCguNAjwVVDDOcvgipRzYR5r9
vl+rAgDNXoOSWKxDnfC4ntUkbd97O+mtUqLbObD+eN2JYosyo/K5y3brf2zW7S41L8erJXe1+LW2
dJwUkjT/vUVOEokngcgA1TrCVWbmAgkhBsE4S2paW/Gj0wrHhAXAFspcCotiuN8YmRhesA3j8Oaq
I+nzr0ZwafxvdbrKmW0TmEZkLpTnbXWBgnKjbVOuyLwK34ZSFIw8ubvlJe3ULt1XbbL19FGdNokg
c52v2Tf18jSnrXj9/qBqFkqCShzVzDGCAXjRFBW+nNNHfQvmLmTEc7F36yItNEGSH5kpi4JbS3a3
XbKXZ+wBKQaLg5kybZ4eTpNEO1+Hadm+VQsCjuDg7zrXcqoo7bCIpVvk2H4vkhGm7H3N7IixFAz2
VXhY2DGAvewY9sutRK6AkzbilpMYGkmY+026XC3+UUsUIIf651N/oKUxGh8iTJVORB9KljmP/GM+
2hVO0Ir2wsqg++LG02HTQ33ArHY9kmopciCc8WmyaHUafNLIIiuiUbND7NaG+vkn9E8KvL9gUWL7
oFNmD5LihoIuSR+vB9metDh2TMBw14h8XjTeAo23MGGDVlH3uaxl4ekekOyaOy4469mzj39QHuWq
sV3Zu7vNTLufUO7ik8ZXVo5PJppHnJeem/a1LwL6bE1YYMOGtd5b8n31PIWkZMEEVPt6o1sxZsI5
dwlQauLOU1yxFQK0noqDn/AGyRbdYeTHtdECTfvmv/f815bDV0yIzjfTOEgwkX2jRw7LxzfwtQ7v
+DLVQ8r++OikFhJR8d3Tjo032EPqLJwTVzSifkyAsm5Od+9zOTxr3HSetIyNRUlVk1k9T2UpyH0C
slP2hxI/hjvjU0B9NLRuj63Au8vMfFyh5lXBCwCTWJx9QyELk7y0RpCU4vuhGHEn5yj0yp/X3d7O
mWLb1gYYLRxDSfnrZygGy7BBAHFek5+/5JCDdOLhkoaxUZvkkBOPGdvD4aKnGgW/NW8jrEoil2Ra
p9lB5xin2cGFAQ5oC0tGob5R/J3irXbPQuQkB6uEz+OVJcmgWqqXJBMsWU9kBkjEzkJWKm4s54j/
B8+NvG92ilayJ+VD9f9ZR1sSwdDHaqR1TarqLxrynuHODRjse7IwlpztxLkkDbpwaaXoacMjn8nZ
mPQFkctSauf1fZB3YmB7/Vkm6aDvowUk7/xKYI+ZcSUCHgq8yKBFLeiRrOoZVJZbEdg4Ibk9jYlS
l7V+1LJlvlnLMVzMbJG7qB4ZyWZf7fclpzbMh7qz4MHND33Hd3oXY+Sz3l6hXp1GJCvcXIlq0605
zNkGumRobGXonvu6I1/eQ0bpawqOVG2TGeB/O7KM52oUb0VV5suhio0jmDeb5KpYKwuqsXfxhDoB
E0d/a127GP3rK57tRAsPlRwEs2wj91hNkz03mCog63h2HdjhbzwK/7oBx502H1ob1He4OGMoMccz
w65o/XBUVYYB+RzhSvIyaZHvEENBDeKlKQJ1imzwt0DN7b7AtMruSqEHvA6yV8jV3TtYp+O8wya3
WERjvET0OLyEFaaRZsc/Q+Zta5XdBKQqv4KFD2pRcxLTLGz614xYSpIit9YoG9QvCLPvJdUMwG9Z
HMKgT5jzgVWrtV2jaxoGtlS62jtZqHARHfawZOl85NbrF4iVsNmWWCBaDr9P7DLdZl7OtzQJsSZZ
S9yDTWc/l+cqNER2Mmo9yHDOvOWy8fPeU5f82nAL+HxPUtNFyaaXsapWDiKcW6Jya1/UIzSzPelf
iKVdLKs+QJ9dZlqA1gqz7ls18LYamw3l6ABdmLTS1Wu7VgqLlX/PTMhQY+aywBsdhE7w0LRziNVM
KfT6+5jfhMg67zQ6edlcPVPx31TDe4iSqQq5CJPuUyhmwn0Xm//oMCL+38vdHz21FhF3Q1GfEeTl
jjDkLqEo48QlrhZKyJ9docHcxs0wj6qDsusdB6izQczYdb8SjSUkJvKVp80vyUZcA2gI9j7FTmC9
cxJshHSIcjvBdZIukXIDH35T8mMz5bLut/eiPEjl5rElEtaZauclMSrJHNkxximPYyUBc393ANFF
n0V8jqrPQRURbCij6suoDqqoQW3QvvVQ2Qo+TiVTB4+Bc3yq3WzQ+Eq9Ms6jH+pKFgHvD3S81Oe/
uBsKAIByW7a7IiZncyjbyg1FKQMZwQLO6j94vJVovyIR/+400rgnB4uFAep1atFgUQ4GwRvR27sd
yGtJNv7imAe+L892LaVIAWHIInrHZnXOYkuE08ymddDaPmmrSEalP4Hr/f/QIoyOWIIDDIgZnkGl
DIibMcnPFzFDDyFFOJIZaeW6cin1geYT3wrz4WMJZhcWuCOm4tCHtrdUydROkIwTbvqrJozVSt9r
3ouMn7PYr7xR0dsnZBOo3W6Pn97mGyxAtQq//W3srBrpFBrVYIO7uYHpJ9f9H/R8s7uF2tP1hd0D
FJIrgPIPwRVUvwB56sJ4gA5rERMlgHMgGec+wf34SkO30PsBcs/KaQqlFr5E82wIU6oFYEHmZf0p
aJ6bJG9Ef4TS4OdV3DW+UjYiaHe363pgiqJ7Ofiv+EJyDpL8LRRaW2f680N2WvsqGO+Fyd0RI9Bv
j8UIdBlGj88kFtc9rXawT9M0MVHLcmQHcv7RJufBGz/AOY70FnV+61YJp9wk9EO9H7ES2GnJ226k
sBpmAlBP6oNwcUlvh/K/OjLJXsdzMnGlnWOIXwCgJFI0AzQjfsLHQgLh3qm8SSDIBqe2Bq+ac1Ak
62TioWJ9+HR+B4pNvdsXCQ4b/2BbeInPyPG5+/9zqtsL+x1FGRAC0s4JpiGsEgCmCZPPVRpzNC+A
WqdE/QbiBwMgah/dEkDYp9D/Xjk3YcFmpfVRKp70oiaopFIO4WMYOJRLSkrbfirTbAPCc4steAXZ
nz67cBTmsSd153ifmNpB0rE1Jlwtbhuw+vcadXbaMtWOMQ9ee5fTfR6XTy3UyYC1/3N6byx1UM59
iY5dC0eRLv4/PMoaMj4NP1JadkYsG/UJPz/bvELOWt1BTs3zSQfKfs+Y4H+crVK7e7/vvy4UhCeN
9SmoRTls67hBiBbCaGVML7UNIKeP9Jof8Z+plTg/nPQ1REw7tKiRN1gq9lXmq9SoydmUWVyJmWy0
Lq8ExIa+DONVnjQSi65k82gRIidkTOeZfO8jpU3pFTvem2WnR25BzQ/8YxVGsi1k/zj0FRfV2aCF
wCCE7VqrI7D/0sGdAA0BHR1LijBLb696K73kEv0yeCgG9PNjA7MACuqr6RE0ldY+9a87cIzv57v9
PhewsFNyxi/yic2mGs/NEKUtAJYMjJNWSUhAZS4DUsa5ztac+Nh4O2wNsecH5+i7qFSxdftA9Nxm
TrammPGWJKbzoFqNN8zLPs0ayZVZWEwjjLLUIXa0XnbTTP8BQkIB59n4VBCKJidcp3yv/aUHP8cA
Ly1caQcYBNZmxPt/6S+I/M8T3KxeRkdHeu7HMB190W06aV1ZK3miyxmjOrPWn+eoZaVlmKDbANpt
HH3n7GyZwfTFgqj6Nb+gXU0rYiR9QiB3tnuRwohDq2G8pIyGB6AEkPogmQzVDq1xDBnl/urIYbA+
QP2QuyO6paxCBbnn/vmtWBubvDTL0OQkVfSHpxvN66kNlKBKugEhAk0znJONB9Viqc2IVsBFPVdy
Qc0scuNmZSwF+xyx+qsQXE6lFshM6IQm6s+DwWn0rvdNJpGtXSHmE7HeoT4tgqNzGgMbxhnppWkN
B73r3tx5v5bzf3caFuTUs7Gsv4uvqnPQHnZ9GHMe7ANKNe2itmqbP71OB5VCLbJmRgIzM1gf3Twa
S1l6+q1u58WXwkmlBsWVYN/sAg/B5ZRoglMUVm8rZ7CBxPQ3ymNEUJ5SKWhFMBnrfldypYo+AGWB
aqZzFni4mn1ixXe93qYfcIBbH5WtrZ9HV1lrGEd7IgZJ7NJctOAEy0tvA92M3RPZdqYZL5XFvn55
VoHGjCWkUV9iZx/Yq2ldlrPBechkJapSDg4pV8LZHs1c3eqz14m4CQo3SllIp+iIcJB7Y2dau7+y
JH6GLx9KBdNbw468vdnSHrh4pmb5yLf20E9NMnanb5vKKUra1lkyv3rMaUn9G9StwS/rvXWTRUR5
1UKJQYvVJVAW7dhNi0ZMdBZAIdrQjZtsYvXgLITuh3YrwSfDWi0qluAvzrbp5kZDSqCM7o+1DmoN
bhl3qoJ1/Up+U51JmuefTdMCaJzKNhZvgr7KkHH9SN1vc3Hq/+uPu2LQ0DeInn/ZZGYRYEWyqh7w
pe4+3/7bES75eW3Kwq2LdfWy9A6sGa2Q0G5PpmGnO7Wi2grCsl1oFRh7KwEZU4pCNKGqfY57jRix
930rnrEZBCbgclXOspKua30Sf6qDr7WhqO9q/8VMGDcMFVbijUrBXDs9jM1O3KYCAu4baqH1uH5X
xcO06IV6vUj2qYGhHugAO7HYFMf2k9nRpBgNVOBHN4gxND7qscvzfmNpVb2aaT8JFO3BTvWQlj+L
ynPpnWpyFFl30xD8fw7togevGE6Ngrnd0XIHTTBCL9EAt1e71zGAQJymuVbzRWHN1m6qg9haFx94
D9c70I9FqPWUzgELZ4zezL8vh+6YcYP+joivVMAHqo5PJppoboXqoiYZVFWc5iCL9xJUljk5jSf4
UvOeerQRoc3wXQ8Wmdx5zgkHwQbR77pWhGd3r/yhMAH3z9P1asvkP5wRVxB6tsZ5zXLt7ODEH6hE
vnd7kIR9qxzEhQVN6wkdezoZw/2ykujDoCsryOZyZUjzaB1CXq6JRxe9LlUjwtIioii++CizEgX9
Qd8IXjBgHWaMDmN+A/DXFGkzgfDI15ZtN8wnxzFtDYbfr5VpzlExX/XsYsNJHkaHs8LVkLAoAR1E
io0rEHX6vTJBNZ1KmSjbP9wPG2E9cMFpLtjKetClsIUwGOSqxeWEqYG44qZKvEhJQwj1NXBx1LpW
x+sGHhFxvu2bblm5zz0LnzOI7qHgZqMC+cJAAOA+lQbH1q6AwxCL1zVuyVnj8+zdtZ93Caa1pBD7
MKxloVgI5uRrLC5ClUjE9WTQgCfIO/Yw0WAznYzKFdq5i7AXgBIqbBEF0n+o5OlDneeP8lUSOd85
uWVx+JxUVJA3GmbhUqO3yYFeQQhWpr5SgvOFchDDKafnl27dPx3unbWp3V+23xVlaGMQB/M5nj2V
dQ+FQilHa7CpBrOK8PBUyoQYLjeGQZ64Z0xzxYAev1iL5wPIJp8cNtnC5lSLj6jFYgM+FidpbZmI
7ccmkk2xbX2TZ8wwvLE7VG8hUiEJJSQ1JcZiFsulqyqXopJlP59lzhI1E66EvAghuFsJ8KoinAWU
HJXzpManEGIXYgefgOR7AB41q8wkahNOjq8BXVdlXYgmN3XP+T1fNHwWQN075aZhKXkTz7amoYVJ
FDnKFCGvT9kgGy8pQrZoOj2BAuz8pCmJLDh0RYg5F84bqUcdw7llLx3m/OlAhe/ZmeIQbqzGKCRc
F9I7l1NYUNO8pJreyUAe7DhQ2/4gykmG+XrVBOyl2iOjbNUiMX/rwaXQZNK6F9ZXpBRdnKNsKQ/2
3O4t/D65NvYtleaN/zCDVvYcuZJHfiK3zs9uOVuoXJK8hPbS2akPcBnX2bdjguEDGUXGt+awktPy
FOSgJkWLLI5Rwat2tkSb9iwrqvxLJAIvN797SEo67y8wuAMdfslajNXyDW9OlJV+Jzsuqt1ha6XD
7bshxulP4fRhXZgFvGtPHGCSGn4RfXY34jPeKmJ41m+PJPrTyaJv9HixKvSHz1uucFlg4w4l/7yJ
9CuRIbGJyZzeT5Gyd7SWWRRmMIU29sPYlQY8ij0DU6+KNXZGi1luqwy1hfry8d2506PHfvFaCubw
8nsjqhH1AsDFiatOOiWfbu+VqVGSnCh2Isb5OAIIiK43DwYadFlGNbZhAqou5iAtOuTbQrqp2biU
TiYyixlgluZJxvJy0dAFHuRby0K2WtatdiSIxC5LH3wlui4UfMHOHDzdrW9LZ5JLV0+OltCgDh87
8IvmBTMjHqwMWwxQu0HZg4aMsHJ//4lyjapyiAQLiV8p9Y1eFPyYbwiNA4uIl2+a2RR2aB0ZUWOx
jORsHxCHK5z+tFsnh1UYEG25EKR2mYfzFSl39BbUOE+TggC7xZg/8Rhhr30YKEv6t8sweJ0f3AwN
PLimOrjFYjzYWYKSCpXu5cGKFe/GL+IeXBuUhiB6/mz3ZbW/s9mH6fl1mKfCqdCxsL39+DvooQUX
kUbox9RPuAT1CSLk2qhJHnmavJHBnZGU9ymZWlMTKFxyBzYtgLuCDOg85PC3rB956cyB5c5htDq4
OJ9CvMF8LyHgFDwYXMvktOoUWXTKVzbH/Lpd6NZqGNwufU41tK/HiyEUiQUiz+chnG5Biqa9RLi5
dbdjz6OwXPS5FE+HY6d6Q7TsD0iC3oCtYooFOyyyk9zDMCp6BOnxeg0+T2EZUoL+ilViQIbUAhNy
xZBrHEstexidbX8JYCs6IpxPdu06u3vOnQPHvSyqbZxkooQtdoBar4zT8GngZTioGpC5HfJS5VfP
Dhn2KCHbFd3s7zN0WD8fUQKS3lqxLFaP3wSrzegbDbnr1XUMou4CezCFkbj4CVI86KLHymTcUfoO
CuXwloA87v4PSgr8FuUMu0n3RKMuFMoFuooMAykC77z/UnURTXOubLc72SXCaOU7jqCPyyqAUIW+
6QClM6nqlbzlEYT63+++OpfUtIZUfPRLU2OZGeFBh7+ybQR5ihGue3oulmnE4ULyJT2DO+SXOQ2G
Df79Obfr6jdJ25mBZsBDhIsRvXaGLiESg1fxSa3F1TWbTs1RgbI/JGrRq3hyonxnS3JDbFyI39DW
UULoaAo6tVc5xKNMpeO18tnx8yiZ7Ch+1gOWqwknzQPpmeu7S6qI3u5hdKuoGyiuW8WWZiOsUKyf
6pGFa5QYlE8yn9oH1OlCNv89iV/1S3ckqI3WjOr302M3FNjGRaioAQ6X3bK0Wn0gsF52NPg9oMuX
LFgbfdWQ3Cd7QylWF0aawwo9PXvvObdT1IEuRLcbNoF2jMKbAnZGMdH1ynZ4XW+T6STycPGcDEiZ
h+lmId21QXOmcxeRUoE8aCkVre5zNf2WvyJ/iLTWU8ykvAxPJ6jcZG0QZ1x8cB4EPZiMekFYNCJC
vKQFhKAqz1xDONfTiaVaBQsdh5G/a2m60owpcllsyivzoiI8+ZqZ1bkFiNhM1t/9oDHRLQ2PmRbf
MYuptXFKvod7v4S1A73blxA8r+B5mZQg5FoE4zSJgOsi8dv/sa06egixk14OnkIvWtoEZysAUhN2
7KJ1YZdurKPT4JcyoYTUjcc1idDO4N8AYC1SZLPnhaPxb3UbXo+fnzvbPv7fpJd8Vb04SbBYGfd+
DzqyCnPyrFf7APhnE1cMw1RbccvlVz1NuFchjYqAsfkW1mhHCINXF+t1tI2IF97mq5aHc31Xh8lm
xBfRptcDkTZ3xw5yQRfEcj5WEao7xhb6cjWkj9gf1oQEiLQBhO82MBxN6NpMCT30uBKsw8Yy/v9v
CWFsvIO34UgtyDVDmL+lTFwGTVOECFwMh4pCyr9xv9T3HQtTJCv9v/r+7XUQXyGyKh4Zf2BO3veK
7haxumCbKV9OgEJvd+Ph9br1XzbaN2J7YFDWMKYKs3jLQZ64fuZEswgwDkysCLs1rMZl3ve0y6gG
qArVJkWFft6Vu3WFonGKJOI15P1fm1umJ3Uhojc8CWaiH4U6z+5U7VJSF0ircfYoSwcagtxEszOE
ihoEF9EScQO8lIJ2mHPCoaTHdlY4IPWjBWQ516GovlQe/FexLkxvZzUtIJJigm5T3+Dt8Pi6SN41
rxjKK0Utjk2IL9/Ui4aTbecug8BWF/Ewac+oig+ut53K9nhLbfW6Sc5Rh2NU+jrGrJtXqNaLOLaB
BUg+2GOiPXn/x6z2xlIiPw5nawLYYlKlAdYzUFZdO1YVV6k81B86/Y4DQHuvZ+/dQAc4XfOOcWhG
gMPJc4OjgsOTEmmpBhQ/53uEak3HelKEsztoFxbv5cqrlKR1vISu4sMK3GxA2lIjfIb7g4IjslhZ
459UIapO/a9OOvdFG9b6mx/pWzi4P90M5xUtpNhYyYs2yBq75b/ovlu8XmTKPI3O3+DwfES2AIK0
b9ZlleyOHVJ7ikU/0Pusu62RHnOUqdDbB/Vf5IyDjteHyVTc21bUIno4AhP0rynAPzeB4enD1i6N
WIajDlhu6dDl8Vyvn3NttsOcxBJ/wnyDeWTuseVh25449lrESUQZvhEZMsNbSNV509MtuS4Hgg4u
MWAiwhk2Y/KkGmhb17iIx2ZSvdxbniWVBM67qdGiJsb3VbkKPDlxeajBhSVGh6JGZ2XcRCf0dlzK
4/v8kagNiDLN/G5YBxKtNPhcYQfdsqasUU/dGH9Tb844J1V3ED353BxM2UsFezDUK0Mz+nITYE3J
4HOyozl45AXp7apKRxazkTI+Cwc0/0OSKPXcilzPzj/Si4mqzpuB+DDpPCGD8/XztObRctZ9QDUo
HHcB4nIwUzKls6WlVYuwkOLW4LDy4TkE2hbvS7UZCUDOxqIYLcP0gr2V9hUUd0n7OGoQyNFGEl4l
H83kCPL+v8aTPMPBYr/rgqTTWvB2LnZfYuNxqmlG5WwgXIocVTYobfqW3Ym2rCxEcP6ibKf8P+sz
gdQZNu+FM6k95wwQ8bXpM2OewfNbO47ke29AMCnqhvYGAcpfdQf4Q2cMW5stdRmwVZhEMqEwegEc
LEdcPy3ziKuAj4kPPZoAvfq4DPrJYEQ1EH7v1Kgqj5ZU1CMhxS+dmZ0nQkSKv4vdc2AaFevAQ932
92GER+nq5kdLkBtHupKzOm8nNojLGNGxa+OFUCf2UoWHmmZjiW0jynqYX8eA6s5ITNQBPI6AHIXg
I/kfMz7Zp1oAvmwHwyKrqlB/nAAhUjBBVX9EPIz6Zj2l77NUlt26P4uje28EY0vjRXQSimXYeFDZ
J4VG3lPbZO2FEVk//TEFOsEP7fIHzWZOb2i480/I7CZSCGQH6dHtwXiHpWihejaNc2/Z4HIjSXnn
mmunP1qwxwmARjdC0PgBzjeiUFWux/yvKPNVJzO71jkEWhJFPTuLRB05aoSKmLPKpFgzIAmqwXJs
Sgx8dMFJVe2HMlHokNmH4IJ9K2ZXrsp4v/kzoUnerbWl4CdN4n46CWR8l1d/trn6CYkU0wy93Zcm
tYmJOIOfwZEAoTdEAk4CvDW6hYPc88Jz2/MfOUybIDY8C2E65se9do0+ahRhx34ig6sVFm2Fr5qt
6fp1qp7WyU4at72EwlidvTGrwPTdyLutad7rJBk1SlvOH2xQ8z7GbnzhjIT1b1GXQYtvPrYhdMFz
4gkZH3xSnk149vs6lunMAgCuDsGJogmpgnZhUe2xD/XnfH8ZRV38CdmzLgQr95NEH9H27j/1rBsz
kAIi/a8IEr5SkEc6++UyEQu3X7aMBO0FOHFGLOaVLM2TBTZRGYkvyeNTrbyIVuASQg9mZwzWtQAr
1a+Dd/7BkszCBUE1H/FYK6uwjrAqXi27YckfdEUH80HQOQzJ9NjMB+6AC0Otbj3r/HSidrost3lS
sgQViri3BBeg/yTDZvg1AEsF5B6VDYk2fuEo20df04U4Qq+AN54ko4JdqmFaLvUi8ApXS20VAZcs
mNzs2Od7zIeZeko9JO9yta4XIqjtJx/QEjiDrtkXcBS8hWVDBUgJYj/1qt3BR7eTqHTprZ6y3OE4
XkKpUXBJL8yd39MjqQDpQXpfg+UE7wj4ViTes28GFuK7OU11Jdgmi6yt6tkMNSBCFvmJ8ERrfvHv
77Id2HXnV/OtciIrs9+YCuGDrvmBzzXrdcEbPzWdJYqUhdMZVcRnkFd6CWrGc0EBa2DabKCI6Qrf
2UVkiA5bSCCC3XkxPD001zYYpHuIumq7KffM3lksaSrd7+jYm8KwAAkzD7HJQbiq5PncXUCpZsVX
g0nKD91mvKQ2f1wrvxOsUKHQS257loHi75xdTpnfifXmhfrb9qvOEzD2pxGQYpZOVFqEbSQh92oZ
owXKwzitdw+rNya4vyZwhpa3+QkwvDVDhH+MURExQMYB64FvNodVOxaPPfXgE6wLzuWEu+K7cwdm
UGgDIE8B08DUbgqIMDUk37bSQYvESIgjyyRyz7HvKmMfl5KpMqE5N4w1arY3q25OV4I2ux9yw5ms
sfU/oJWC57S4jseHJnAe6iqur2Y8F/XCbkLYvKk28GbW7N3em7ki0tiQIGGdqnIvbxpWY9zupdSj
IoeG4FaUVKPwBicNmqHqhHdfoL/LNk1e03iImv0ykM5fD4VAAvhi98ZRdHyLOxdcEK24YVfVHLVx
2nZp660EJ1ZZdDZKa+CUsYyl7Iuv+Sas49/5aNWYaTALurGEuimsPgdgNgRYIRpd5SRxKELJs7oK
unnefMeUXncWyuA3pvE5h5myU0pwkakWinJx0gSyIamr2qoe03a2lOY/Muy6V5aDCMk6ekTlrAh6
TTCgzfUwA70Hijt12bbm8SY4mvG21MjBPcli9cPCcujyMZU/3nmxZKvVuvQYcOnMjj6s+4l33OHa
1y+GEHpGrNtchmEVnJs9d3SW7oCaDvGR7legy14SR4a0wkIyGNkp+Jm8rCWZWAZfkL0iVlyFgEXH
6xVey/HR0djUF7MhQcVK3K8yLu08IFMpxVlmbrx1nWGuYYS15mHbRF482gVuqgSiMIo6jV/bZBUG
7pMLwdbOQWeww122N/DRDd66rQUAjJ/dhsE421DhZt/S77jJtiO0pyyBpeY6UhERdSBkm/inW1TA
2m71b25PvccK70aB3x+SrX5PwJU8wn4Q7uX334VfHFqeP6sR2skHQUE1FGzw5PN1Zi8Fr7SHeDgW
Q7bnUx9Dh94CrNhcMRFq0vipdc0dKKAczYC/v2eX+hqQalKt/GkP0PqGaCb/bRB7rBIwm4m00u92
WzUmy+a7mm3EMDxjhrQXU5B0BjXonicKtydwe1LMhgOZ77AKERNKDQZIpCBiUNnxwYT01zUSPrRF
3MLxqFi3QbU0EDT92oCjfc28Mpl+PZtyM+Ie5oOa/f22SktBkmFnyqfXIRgvOCzaGj9Tz+qfG+0y
Zr9SLzhZBHpt2j/Yqz5Bf3CJeDEO6eil7lwfQaAv3rqoIF3oNauBLzEzAmubNw5gW8cBCLGyKKUZ
lXW5Bv3dG6IC9ush6O4sDIO6q1N3+fOq1TWxZKy1tkLPfyMPIb1C+DlWStZIktzIC37Vo3b7cjvQ
9/vvOUBCZe0wZrnOD/YO39a143YsgY+N4Kd2ZPRnShsm93FzmuV/2Z2HSQqfEyZdc6sN9Sm97Ug9
fgHne81aIXWz9i3v0d7HXmS80nP2bjxpFaaYWZiQKJmHtjs4s/12GrxHiHZrOQBkniPF3CYvjK+9
zveqLdFklSnP8ICGUsukQOODXyuIW1eyW1Xm1JHoGVyySmiGk2sb3m2qCVTT1AMnbrljguEjt2ZP
l1taD5Sg8eDeu8+OsrhVlCxQOisIRF2nUV1HNUjXv6VXhHU3nOkfEIzPL2WXZP28ZxfThhyBId7C
i5RhlHCmy08r2lTSITJv/bsb08BSulsOPjVG/rSpzmPJTIr2pDqFK7DZaJBchJDoJzTRWDmEQyCg
fWbMriikrjP59yCq8w0+6u9X1wd+yFVLOULnZnvNYVFbnJjUUIhHebHNd+W9pZ3+VyNSADIgQodG
oMc74CnrQWJu0QXD3yixmk459SxTmdE+EAoN9+QwYKN2dfP6MnOIo02D91hIAPhJiHcT/u2FbDo2
7JX4DM6H8d2IdllyIsd1rcRUDgdDGQlYPgMSDIgrLGIzZ01cXjtExbD4iw6irEmVqWLyeb1armYf
3FB6FmX8CCPxWY/SapQeO/Ibs9jbhQsCJARuEJyuDjr48Dr/CVOjlNM0DtL6bQ2fzpXvDX2ixw3Y
SOKAG1D0DaY7PkWTTa3q+2nfmmg9GAJ86h5lQuQ/EwpixRCZGesXlbMW908BoKTSzSuM8YSWVwel
YR8pF98o8ZYL3GJBDx6ZM69ePJFCLZmV96vO4Iy1q7LZ7VhGNkBcx5eFDJj5u/MWMyQSAhdz5OJv
HnW7+zjp0GWF2pAHna3vARuEZ17tjf5/SoEVNnyDf54er6lhZu6E5JBXbz8xqg7J7KCWuMTq/5Fd
0Y8mF0HRS/VYhxvPPKNAjFIfmStiIvy+n5eRryjNlaYz1WoqKz354j6X5PD2vXwZamlnGquSQ/Hh
1gxdFwL6LyheEO9dT5/LYakq/zluiyKqlC9XacUYS0UTJC2lYzOWnHzlRlyodQ6GXDu/ib1lG+dl
PwRWSX9HJDW57+aEj55X6aRC1tr9XVPvT2abMbWsilt9MpgZSN2YTczueEO9ou2b2f1PMXmz05xf
S28l5j0wi5y060h9zlWTUiYnq9g5QR1DHsdQZRRnuQ0Y3cpBdUFaPu1l2H8T72QiDjJwV0G7OfU5
GbMIvURxAdCY5P+LSxirZ7IbBF8piyIcMx7fWPO2sb52bQB1hxHr5eAbSOoNgWgkbWZBv1QSRBYs
P2OzGTbr4Avlr1xaEzXw+UGWqT9X6PmPS+TIzgBKo6CNc+gVCwEAI7bR2oib5GP/NeVyb7gsPCMw
YBoe6+bucO8RbRQmTCInh17A0HIJPCgZ+E7hs26YUtnYlfaK0Bvzjdkce/tUpBlwaUEz/Jab0l1c
ofkpygMvNv7eaYfVIu/NaHFRRxkvF+uJC7VIe8/wtt8arT22m/uXiFw81494njhqfdLk6vu1dgrk
ND3DbvgfWZEJpOVjk6ql9n+f+VarRLWvIgPFXckdvXB1vhoGmlGld/sZIk0AsxG6rFNDgl4Gnbc7
D86/h+/I1Yw2x2zoMCPCVRB0LQfmFNqf6oEguDjidHPIU7DD1hl3P4AOckZkPr35dGNwYcJoCl7/
l7A5jgVDNBqHSm7bfZhVV63nCtJfkXd66u+AALCZ1Tug+FGrZUHo3RoxUZHjurt6XSSMv04P9Zzv
bg4QME65Cn5d+dpZFUFmFfySjbY1g6WrHr0T2DeHNS5FCHUmUzKKMqV6pASR5uWemH1ugsAU2VuS
NW7DEkWQPTwOLtvpr5z/hBfgy+TI7wb/+R8xeR/KkdJ3/0p4Bz9uktOjaCa/cv5xJkdTpzkraOBk
ArjHKD9ybiT7CdSvnX7udxjt46XaJ9JzASe6qBiOhAx7dlgzqf3LQjWnIpiVT+fQVDXuYJlkr60s
vkPor/tVEmxk42/9xLG11WWuJTgYpjBSZvcYCiO+qCxGVY6lIdBl7QZ7MC4V8dihs/Noj6rZ6ApD
WWe4TgxCuXcagQCkAWSaSN1yoIqQ0uarh2eDZPxZSd4r4Ew9KeprtThDNCT9KDnC/eZMhCuUo006
hceEk4+jFvhEV3OHRNgaDGCXQnaxSjzw9z5JfENKZqfNdi/fuG/dxGBOWpRVrcYDxo9X5ziBPGBb
Ck+746X2XVy80+1t5Rg8xuiJLiV28JFmIqMYI6UKJuTkadZbU+AzAgjdQq9gMkPyCo2gAFTZ6y1G
HcRRGlfI3kiYF0xnQClaD53puOSPTMX5s10M/YiaWfQdsXUKvwQNlaaM4svLyzQ1dMJ0fnLyGhWe
4q+osSy7vKEyN2zdKh/SjIaouHobR4FL3UI5Jo3MCDiu6ONnbN4HeQoDawE3QuyD25fmC43TcMfD
87dDZ4QFAQeKC3cB3pYtl5oEtQ46fuVgGjcl5Fe2pkNKczk5A5X14k4168hq1Y2b9M0CkzCzQ3np
TECCtvynVXzmiX8WXlLHRa65Z8hExcr9722BqctP6Ppd2OiwMIcUcVbeTekpCV4kJjuFua5yOh9R
LQ9OBjQ4JzMJ/g4oos97S5lNQGNsttxqHiJbkQ8A8K40usDXXkrdUyIW756hObPfobUaTG0bkbkz
8n7PlzRxu6u3z/B6LYZ8lFgVABNd3V5P5ELvM5b7yP8BCZ5G9E6cKSPE8mLIgOajLsfl4OkqeqhE
3RZDIcaMCweFK5rr6QwLNB/lLrAl8eIAzFmrAm9OxJavaD2m2n7ZBdaqVcH6uqrzx3MmJ2CKhDd4
IFmhDXhB5tn41p3qnjXu04HcDxUJizpIDBnXEp4JMTawFcMMAAa61uKY3IJ+FEjaTThGJXviD1Y5
2V5IVvqY95FV5AGbaqCeTIRtYT6qbaTUuBE+p5goyXK1IyqMDx3wdXdowC54T/QmBT7po5PaOTVX
iGo2rdMv7D9OXbtbWerDzeW3XuaXyFhShFGTVcxWnaosxXsm26VIV25xkyGEUDyIs2Qm6uF+GK2k
nlzUmDfJnDrBYTFD3OtUBJw5H5zpFEAeovWb4VlafAXshngnAcQE/ZNIlQbkdLwv8le1lZtd5Msa
tReBUpp8TRHYQakauOyW3YAjjUdSvSwqdU8vGIZ26J+dHvmlBVuI5fLN4AAQ2wXTB9gqWpwBpSwn
EvjvH8XonCofy42n9Ej4jRhFXxCzuLqx4fQVayVkyTR/puLNfqhERAIzFCFvxVPilmtqvpdYp6p2
XEGN/sWrdwbFDMe+1ohu/AvhxTn7JH+8HCBr6xejCeT08n7UMuY5gstCENGodwWoZznYmUu6niJk
Jb25urJaRTPDc7biQ6iOl/xhRosARCuFQz5cm7oTHGQNIYxqYlk7vSnc/AiVouI86IKBmFmPILin
61jdQ3c23FU1XOY8D5B4CQeMg+uAnYfKYoP52zz7aYCdrOXq78MAOFNnzH5qcXZCHV32pVhXDLPF
BuM1iktF8tUG2Rj2rRITs2tChte60PQEZ9SXz08IaFX7G99MqBbdLJulsHKow3mxiPHDzFeSZ1Le
Va1EnfTpGO+xUugMimS6YoqYjP5LsLFsbEFxOcxEoKDtGZorKH1/23O7K/dc9HGd30K+Oq3qlHi9
u8mjfiNhecwlERfF8flMEpbJ6hUwt6magODnb7hTJLA0tY7Zd5EsT+tMgd3NH4+IHbjfIC51d5a3
7/Wp1wSp8k8ZN57gN2tYaQZDxqOKELCngYKWOBzerfWDvZg5eSKi+dfLTaBQfvk5X+FwDhKtZDVu
Qs7NocO7j0e59yYTkOZyQw1JI60x5b8Vjixe6aXYrHWk02xLDxu/AqJqS3FeW1WIXBEmZYGRMtJJ
1kN2Wd2v9bUZeR2YgHmaHb5g5KIRf0+Qvracn2iJ7IHV4bxH0gMGFiZpKf2ujUVAEx51T8LSxyny
ECN9X3XPIACtyYZX0vHLUhY88Z8Jy31R1OdXNxrLeG5hi5zPzPl6yAXpSifJQBtuz7HSkCWueV0p
YsPy038EDt72kdsgy91D82V5a4pinwyUcV/Pd3p+IBaZBYpbE27yKNoWr5z2po6Iu9YOrYYcHlgh
3dPhnV/Vez7OcVZKRrFn2sE8Tyzq3CsF/zFLejPzgcFYdMPNbR3QL5gowTDberixjoIfLxv+pSG4
+TFZRZpEoJQIYBobLRewN5tdomQYcCDrvk/6teRDgFh8hZA6D6+VMQcJG+62kK6bGbdN0A3fnyhL
qZ8IZXq4s0fRl7UzOUtgkzH02J8/cUR9EkkN6z/qlOYJnttGzLuuTXUiDSswLHrFR5AgXo5YEBo3
aSZidncZjGPqHhbmpAom/i92xIdQyTx1LZrO+r8bKlyMzjYQmHS36/6/fivBEdXp0ppraSZKEhqr
M2V7jcdjY0nEBjhLkJgXDIi5zpADMYX71/wRJzEXkkRfSMWxuBdnFSzYWlc7H2W3FtwNyn1cMYwW
HBAL9hy+Yd4CCPGfp2oHNXQbSdTIzpe3y/UBhcuSwswsxJefOAogHc83f0kmg66Z20IcD/Eh3ECl
LgF8w3RGGk51qWy/gowSeXwkYJQJBOB0XgbN5AnwdcZlPDL+aUpNLEwlb36K8SJDbK2D94Nb7CQQ
hjUREXkQnwyWlJNIHUSRV2HeIp1hX1iXJ/zlQevx9Jp4OrEAYm0kl91zc/3yYw1aL0/MDz6BYbiK
1qKHC7/FZr1EKKzv+s0+R81tpinFp+YmoRiNVRpGfqGVuApeIRYNxjqnJIt9rkGleBvF0jNohcJT
sB7jX4DE7zulVfaLAVHUr7LUv6bRYq3Q8pehyX34nPaUorrENEBGJnHYnYktNc5JfDNbEqZyOJkk
/W7h7mm5IQdB5vI8z6IFpslGcX0mE5lcMVUfXvE1tl7XrpXnyW9rPsgXNDAwd222dB2gZd4Z8Cz9
JtPxqc07uujPTF6h4d96Zl8PohONEBcCwmUczj8H06Uz7bayo/0fyKP7BP6/CFD0pZfEZtdgiZfj
D7nxMHIOnl+sMfRt3kpkJwMMW+NekucT3o98EkbsCWTZ3bMAm3RTf3TjVyBrlWZE8EaOLEAIj/8D
s6DOPjGtGSErujhzzCArNYb4TgYq38FJInWr7Hg1iTwLNWBe8LyMxMVODqJJKp8RWhiYzPsLJ3ae
gUTrXsPixgVKqTX68ECy0ffGuQK4c7rUih+c8/+K6QUWafYEaQ6Tzmx4ufPd/zFxHWsSGPw37989
qmlUEBWCq5b2jeI/07y8t+J8d7E9VkZzbUIJvaHe/f7IVP9aP2r7W2d56D+H912gf4/HzqBrn7Pf
Wql36r6aONFlMJkgHpcLbUdNJHkJtQm8L7je1D6LDGOq96XEqvnpkGiLx9OzdMWd6Hj1DOK/zF8L
i3a0q3mWDvQjmYUvY4I1Cvgi6W1V92eXq/5S103VTS1gOL83MsvyPwTVJs4vgx7y+YonINHaDG9b
qXd7ZU7f4GGbu38bepWvM6SDhRbVvEYJm+w/l/WR0OmEqdQ6+GZywWmHnrf3hUzC3Mhq6a6kOwRj
FQpOfp3ly5IOn6XYDcIIhir/kvHoqpeXgC2N0UjrcVfE/kOWY3pmaQlu+DCgVClikHDKZdePDaJr
aIflk9vUzX9TmQ54RY5c/PR24dX62p+3vsvF7i5pAS2nC63t4BXbE4EvQ9FM3cXIQjqwD8hYJNpx
nMJNHLVivbV1/lTq9W2ksIWoIoAjWKs11IW7J252TyjEshcRMGGyDojBn7bV6GUxwmG325HJWI3m
yiXXLwezD6gimb5dbk5uVMe4pjKgPFSOA8TU+f6fiQO+jdSxIzt9GyJuEk+mbPgxf0gqUUA5NKYT
DVZBYIsw96epvG7/6NG6YN4vUGQr+8wrVaTAS+nfg14/zr+cKlTnzDZdoUcEWn6QgWFEHFwvypek
z315k5JcixM9CtdKVME0Ye9heZyHKUepLwP9pr4lkmjwNiR3aIAvbIZuF3dtQatZeOn5UIAqIHzm
i/aoxYVWLrBDBvUVCDM+CA8gonnRkrVwxbI4nN54PEhclzV4tP4xl5RNO5xr9EncgLFkMQllmFDw
FOBLaaH3Sfc+bWp8mRA5zfhtn/DPGKQ62Pj+o87T+B3G1FHlDV+023Dp5eAvRTAmrV+xNN7+m2Uy
kVWTppjehSfZCtD5iVw8TQlmfXyW6c3yGMARYm5xlmgRwEv4cQGkPZCQHNO+ICgEr5YMdlN3IUqc
YgfnMOtji9SAI8Uy6G1Cu3EiC3nSwrX1i1U9CY4W58y5PZb3sLy8nq0981BM79IJJYWrpfqm4OKM
0vgYAFAVvq2lSE1t3qwA64WyW+5GXuRD1v1DPGOuc2UJF97/CGh3uOVSnfiT393AAB6V+uCpD+OQ
dpzTEL6oRe2te/NeDuUCBURDfgrNG9/ndRf8rd2l369vqo8favWMhRA7SDKsizgZimymwWFHYRFj
jN2+gu4bWAxi/A2kzsyWPfnpEE43OEHXWRDm3igdnYkSIciQjTVoQygLZc4xoqKqbY8oarV5CYT6
qtFBOdoGQBPRq86Dr6eJ9sOX0jj8yLhKDWqEHDq6jmBkzB/vulReQoEfaJAnZ6dKmpCnbFpt/RKF
1NuwLTsnARFab7wSfhlGsUcha49dfKuYF9taOAFrZ7c2X5tmH7p4LJYmMvwoERBSC+qQG7gDpmiE
MmEBCRIjqjyo+VJfdpsbnaNWvLT1ndRPD+Wskjo+UkdNbFIQipbsFWrmrPChK1IdRm5s7uyvzzc6
cgnE6gtm1/zKZHxXMRUudLNanYJlitQv/qqspo5ykjgs+vIevHivvt/gH5m4+hPaEZRDWikswoPY
hPrL36cRS0W3Ia6egDShNyLlSGCPPFSfkCF/+02n+KdkghcCcLilVJSGLSMsnrwTlyqbfa0gZapt
1QVZyPntrJ55L5zlqtXGzXh+Z3+T+dCiE6cAdRC87I46wIM+jLkLwmTeOtT02Z4yj7JGkBs7DUJY
EGaDuAbm20p9g+s9K1TEPfkIJOjGqCu6wNeLJOdUZCXRat6ykgaR9Ot6QZXZFcLedYCYicFAd32b
ljSLjeizn4fmP1G5zY3xtwL/LrUVfXn6AZDVcOb7gH+FqE3jrbDWJCc66CsLN5hjVZtZp1BzasE+
bn2jqmLbKeQOr1bSZg9T/jvAmmHKFP+W1J+3V04nRxNZGG4IIAg33nlW89udBuM+NgUSxGuoYYjD
gpZoOBuIwHNzgZqzrerzeY38/95+2l8p5iwR7ALE9/y0rWpOvEdJxXcHSwk0/oHEskfkBMxFL0yo
qog659A6QVto6lHPzhYCS9VtTRJOR8/dvjKuUtSXh6FtYUr6JqLNyRMP1wyvbKr+vf6YL2W7uvNC
FMc5TG752QC7BX4bqVf80sFLaz3vb5IudevIIVbRp/f2I3K8b/wu+Y9cX6CHKcCdQ/VNeXEfjpqd
BlyxuHmkgQaS92dUwPqYSn5nwQ3ltWMBDVAjhCp1hKW7xAa34GCmjuWdssk+ZmXM0FcG0VDiZhyv
JJGA0vBDdaMn31h7Gb8iS2jssrTGHPvAHn08FcG/eV/OlzAazQncN/+hTyl5dy3z1D+o3BFomkzx
07QbsHBMAEtlc8RB5Y7vgIrMhfeHGwpkonMnSIXItaOyWt8Zeqpzxyif0u3dA7ICMM8QJvNyaeCD
upgXb2Ay6m8Z5WtgnBPBobUyEQGqSskD7nePpC/hk7+7KdZLX7wYOMDBOQF90GaoANfPHjYednoe
5fvN1vomGku4QAziUhCIQ1CS39eHc9ZE5MwpZ+ts1iva9cN2TYMxND9QNICEpXuaUOjLyHhGziZe
FAdrOW8bGl5oPc+XW3ltDwHii+lKEqXtepcS/bvnOiJ6Kh6CPH9Kqz2TUhWNyBgfm0tRcXwVhVRF
vwGlbOFF1zfMaXyDiWwmkPmyF8O3NOdav/jhorkP5aicuRBKCw78FP8RxjTM8XXRMG1XRDgCIl1M
4vdUoOW7HgaV2e+gq2wOhHeL0CRPTNmOAbIYM7rIOx7k1mNumjSGTp377+FmPsLCW+XLbG72LxRB
yLK7G7vk4DCEjyZl8GaI/L8fu7tn2zJ3syhR4vt+hoU9Fq2HrVbnhztCaBLH93sEwdL9t56W4MkL
RTzsi1BG45QcuMYnAZQOyUiIAWtW4iVpD4kib6iHJvt/hc7rbI3tbYtYMVjx2a5i3okroV5am5pQ
gNMTJ07wvSI7Fp5pwW+fQfOJZMxB9SCEvVyBxoGSWDHJ0fWwwbU/RX4wKaFt1hPWSPsO8zs1ugOv
UexiokK3llcaNYYY0iamGTb7luaJTM9iRbqXcOG0Pm/2y93qwvDcJ4/GXv8x8HLPEVrI0BT8ZNlh
htgOM37adVONg4+JJg9UuwpVpsE9nuJJnP7aUzzLo98ekgbIlsM2oJYyG0jMLydCYwkzY3X25++Z
6mneQU3e9xDZivpfv3/ZfVc7cekSp3wOSkGUNXpg/ij8k5x4lXumlHUfBH4fhIJwUDRtJX3Tb+6T
qwv6TURfrOeRcyesAvnixxfOaeL0ZaTwWl7YNBg/4RwTM8wbcMi8na8LeAdFLModjV2jfv1ysuua
6syer67frb+9hjOX592vX8n29y7649LCXvBKBsOuzJniMdTRCnYjcichfaRt/eBMFQczsSnGZsLE
ReB/QfGrHtmj6dG8CJBY7eIyu0WpVnNbCE5McOlM6ewbuPKqZL/O7YBm4mWF751F9DweRiHcddBB
TbSCtlrcN0Xc1xcJ3TIBkkuFmmbx9fG9Ruj62xKRj3WKD2AFYydgUCiZJ76p8HkIZDeCgnf0pphr
fGWMd7H4twIoCFFwQTkmIDYjFWqsrn6s3Gu1bN54/QZ/CCC3u3AUNgDN0wZfAiATJxMSn3mlj/G3
MdKEQiZeqjLqGvIridkXaAmYPV+2o2z5aYAAjLUjuQrWaOkPcf5zLGCDHp1O3KMTbvGDddK5JeYg
9hj6XuhDyfitzZrZH9GZCbGTjo5T4SQHvwTsTtwyPYtRWzumcQ4ho1UZi34/kSMkeUwYlhLxIhYG
+Nhxn7iL/677w7YNunVANs65kB/z6EaFHGCr4UV8qyBHoYb5NUqrpbVtOgNzTXvtGxRh3LuLF2xJ
C1ITFhXdM3j67CudZyNYWVmY3/p5VezJBGMcU+fv9g0tHiBrndDGX0IysECFzSyIPonjDccXmf7P
HjZwUluoMnTgMMtnJJHJMKYTagi7rFRgVtx3W3NKywzrPDFpY79sYQDhh36z9mj7ow8EQTe7Dm+e
GWd2FMnPS7PojGUTS4a6653pxXyPPjNHuuBToDgL41Db45ColKP6Obx1nzhKNugE95c7050XhR2x
MmivIMz1ALtuetL9CAe7sUYtg8/WgM/G7ZuZBEYhErf4ydA3yMxYpVqzXGVM9xm+sBYFosEYQeH1
hEf2zoaySOYmZKYORQnK9UjAmrvgSDMFK16tzFFeeo5/pe0GIBs0w7FODVAeuL/kKpgfLnqNEZu9
2rZUs+BPKq/k2vgK+k+4TS307jnn7KUhl5m2LY7LaDR2txX+nspkZ6CpLZJ266vlOtthM7s5o5ig
sGLj5NYxA43Vuh1STr3rGOV0/oU8n5tBkR1mKSdlG6OkElmng09ByIwKBJNIFdouHgBTwCF5SsxC
pJKYePWKKw6pUP7BVO+AYP3AXV1BwSCSwHqIXI/IbfGJ+JGgkVjsa0d4ieQTvnv8SWBJ/hQ3S6D6
8UlJS92dRtk+Y7yBR8ksVkNwIMseZl2EY6ZTkCbeRtlK+cUli9Rh2UYBBT2aOXg+2JsXzP2dKUEO
YjUkWbtHTgX8dtdntKLRI1IZ+Ntwwwdi0FkU0WCzHkBox5KNHjZZlZ6A5x8tgiy6Wk449tBWEJMQ
j8eZeAfJA/ELnMAu00P3kUDPXYTxrutdVcuojFAWSWQrC4e55Az1TLkzV288t+q8v04EcpBHv5c3
ja8Rgi+krdEwFJn5aRczuE8BdOZNFSVPYpQ2fDauxSN4g7iJ4GzpoJbAYJnG2Y0m3H3cDH3pLV8P
FrkCHOgACxlajdha/3W80YpTmDyoW+nvDSM1ggJueC5KR/uRFWLa1c4LRtEU8vM5iBTLxN6INWXZ
gA7eOC746flKDljMb0LjcmtfhE04o0pu+JOh6lpVRrhRZORS7nNGxvFVek8EvhEjph04z89yr2MO
oJjU53bPJYdE6a/j9Oxczzw02Qi7sNuRaNO+Q39UZHtY9GI/ipHMouJMUq/exOl+qjxZ3EVF99Hf
Ur+l0fCHTdSriLzYJjriukbGaPI3U3zq2PMZtmq/JEqYQM/DdbtI7tpgMQ0tL1jKZtnyB4ETSlhS
j5+guK8w/H0daT3aptJ8Nr/NkKw31I3YwAJk8ML2Hshg9TmRTdnJxXt/N2EfgZ+/sImJnzhZ4VT9
4VE5wrZRtlCVv/EcbIqtzQRt56m3+5lJefKTq7gN0PCtQBbH8xbRXhrXF12JuEICIQ8+BuPNm4TT
puRY+IGN2o/HHgBe+3YYqfKaFysTdCT8mNMlddak1paqTQLJL4jL0Ks+FwZsUdQueefLG3/aGFDi
i325ND9cm1ReI/Tu9adtKHsK5gAZsqbL/ijtnEbRIv12erwcV3W50tTJRAO1fT5amwZnjBj9NZyC
3dhIuJOGW5xLvkwrtAMB/nPlaCJRrhABC/iBmcwJtjo6z5Czjyl6rncRqHDnuoHdaOxYvYwRwW21
0xTYn+iL26rrI0fSzgd9h1H0DvQ2l8feOprVRwE3jXm2U1FOnvYIFxizsPIlNruOC6UTIszJKMBN
KH7LPe4ht6R6GNEv3K4iWGYZ2W/KZ14YGDCWGA5TL+fkIfGGD0Od7U/u6jfJIvBxg80XBX2LBJfU
06E81iXFUqvy6m5wT7HJ0vzzRS1ssMxF1pq2yjQSnPCWg5n3aNeQpNKQVFnRcp2oAt5IyjULeTEB
YLmx35z9bdShcDmwgKDH9ypj4KrPf2nNcdVKNBQ/QtK2AK5/3PmTdVRJ2QTvODhRkanEpzKQ4ldm
6TVPZxly6ANpSwebRjTrTwoI+Ke4uhITRWfk6o+qs9FarIjALWbzG4wnM3UbuqihTYz7+aaFUef3
kY/H2WS1DbAVUNBDxTLd78wM3eLZ1e/ffyx83P/WcqEIVhYf8cx6PH4tu0xfr8rcEQIIKhi1KK8V
OIsWpwedlSgAPjlNTDL0sWDMKMyJfFHRGveTTS554jI/bFOT++HCYgTE/ZN5opLGH+ibuCK+bJm7
OLnDq2yTzrlCFnS0rmcJOJzKmSglK76akNwGBMYpq9HAu4Cy9X/5/38vCYZ5ooxq3n3lSTI2+dch
2L8rFm8QHhePeg3yl9mzZMTHcSilWYN+5ODOPlYgVJYAWasnHH1aPfIOXTpoYj+X8jKrq+Sqsg7P
vYupEOjYX9T6B2bH7C7XjTrJkf0kqnJu+hojXcv8d4BjNCuTVLi0hV5BxDyJEIYclqVGhbQna1XJ
SmqusPUrY4GAAQsR+88PkUfRqugAFWpIxmoRQvxLuGANsLBfA7u7ImWF/KLeAdxRu0xeEJnH9KpX
jSb2A62mKklWDQKpQVA1XgjcTokwiiWMjYkAjOqIRfxOABu1RePyt+bgtWa6EjhIEpYbAtltHSdw
MfimIIGxsohO5V8XaSLsaBGA8LiDbCINQFGfQsZyqSpHG42mfZWNBOB7eqvPg52fvjySX/6HFQAO
SsLFiD3rcLbrhBbiMF8kTt981tYqSqjwyp+rPYexuED4a6Shw9uJll2hRDZehre58a5RzPPolWB9
DyWFpihO2kpizN9W+5u9OI6/wiNtwoCQYRm0D2g5rxcWidHud1kphWIL/z9ZjKm8SpcNHvMcc2hQ
qanWs+0d41hLEWNVaNxL7OxVNReLH0q17TNMkuenAxsFQAX7AWyneLNeLJ1itkLuqMcqh+JTTS5y
QRlVmwhgt05OEWJnqraexoVKtcLg1YkLdWmZ6M4ej7zaPyhROqE5MTd0oLNxBg8xxcNpN8ncCHDa
hNhjbM3YPLPEHffiMbGFrpGEpyHpr8JrvnZnalFsimeJiqLI0tpYztvr2NwKkjXHYlskuEt17YbD
eoPrd/YJKw9MecID/nwupIkNoMI8zUVSEqXOiXrGqMwDBvKbY11jCWJYVywLPUZnms3QkeAowzMt
EFnjTFw4yjHaDmVqXy0ZyiuNunlcA82QW5SWZuEMHri0Dh0hq1wtbIRnRKUSnvkR3MapP6v3iV/H
zg8Tyl6fgRudc0IK9lrXJ6u3MgGWF5zni82WmOBfdep0l+E1Esk7iIesSd6BlrlE0mW3UEPCw+5U
DhLbtxdrP0I1zaMv2X1+puuJQlFe2kQQWMydFFmMhaBrnxaPH3+8XsomzjRWnLYVS73PjeDsppS5
O3SbhG3XV4nk2iMTpCf85GzUOiDFN8ywcwDiRS2IeSOCZbGNb1H+eJDVzKKIBbE408LXmmAnb417
nMB9aKMAxR8t9Z6876NJyZD+sTDM2AL/kp9PCzTJB+hcNuVd55wVIoZrYKazfDHItRENfIvgpMac
1XFyXcRtKZ4Ty50pJMF7is7oKshGyelYTXiY4ISuShrweM14Xwxv3GKVS/KppgY5NSHuvVyV0mtv
KNWDp3cD0lAgFuO/q9Uck5K/i7k81loU4v1ZJXmd2l/FRS6x79awGp/od7XjHjNvIjzjdbWUi4JE
awQA1OgamanATkCS47SIdolzoTYXfIxClZAKHrRNKSBb9WKFXz++v9QGnA==
`protect end_protected
