module ila_0 (
	input logic clk,
	input logic [255:0] probe0
);

wire tmp_clk = clk;
wire [255:0] tmp_probe0 = probe0;

endmodule
